* NGSPICE file created from tt_asw_1v8_parax.ext - technology: sky130A

.subckt tt_asw_1v8_parax VGND VPWR mod bus ctrl
X0 VPWR.t28 ctrl.t0 a_264_2813.t1 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.5 l=0.15
**devattr s=9900,366 d=18600,724
X1 mod.t20 a_264_2813.t3 bus.t19 VPWR.t24 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X2 bus.t14 a_264_2813.t4 mod.t19 VPWR.t23 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X3 bus.t15 a_264_2813.t5 mod.t18 VPWR.t22 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X4 bus.t16 a_264_2813.t6 mod.t17 VPWR.t21 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X5 bus.t18 a_264_2813.t7 mod.t16 VPWR.t20 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X6 bus.t20 a_264_2813.t8 mod.t15 VPWR.t19 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X7 a_264_2813.t2 ctrl.t1 VPWR.t26 VPWR.t25 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.5 l=0.15
**devattr s=18600,724 d=9900,366
X8 mod.t27 a_680_3582# bus.t25 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X9 mod.t14 a_264_2813.t9 bus.t17 VPWR.t18 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X10 mod.t13 a_264_2813.t10 bus.t0 VPWR.t17 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X11 a_680_3582# a_264_2813.t11 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.15
**devattr s=17400,716 d=17400,716
X12 mod.t12 a_264_2813.t12 bus.t1 VPWR.t16 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=52200,1916 d=26100,958
X13 bus.t27 a_680_3582# mod.t26 VGND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X14 bus.t2 a_264_2813.t13 mod.t11 VPWR.t15 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X15 VPWR.t14 a_264_2813.t14 a_680_3582# VPWR.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.2475 ps=1.83 w=1.5 l=0.15
**devattr s=9900,366 d=18600,724
X16 mod.t10 a_264_2813.t15 bus.t11 VPWR.t12 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X17 mod.t25 a_680_3582# bus.t23 VGND.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X18 mod.t9 a_264_2813.t16 bus.t9 VPWR.t11 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X19 mod.t8 a_264_2813.t17 bus.t10 VPWR.t10 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X20 mod.t24 a_680_3582# bus.t22 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X21 a_264_2813.t0 ctrl.t2 VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.5 l=0.15
**devattr s=17400,716 d=17400,716
X22 bus.t12 a_264_2813.t18 mod.t7 VPWR.t9 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X23 bus.t3 a_264_2813.t19 mod.t6 VPWR.t8 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X24 a_680_3582# a_264_2813.t20 VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.2475 pd=1.83 as=0 ps=0 w=1.5 l=0.15
**devattr s=18600,724 d=9900,366
X25 bus.t4 a_264_2813.t21 mod.t5 VPWR.t5 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X26 mod.t4 a_264_2813.t22 bus.t5 VPWR.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=52200,1916
X27 mod.t3 a_264_2813.t23 bus.t13 VPWR.t3 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X28 bus.t21 a_680_3582# mod.t23 VGND.t4 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X29 bus.t7 a_264_2813.t24 mod.t2 VPWR.t2 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X30 bus.t24 a_680_3582# mod.t22 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=52200,1916 d=26100,958
X31 bus.t26 a_680_3582# mod.t21 VGND.t2 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=52200,1916
X32 mod.t1 a_264_2813.t25 bus.t8 VPWR.t1 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
X33 mod.t0 a_264_2813.t26 bus.t6 VPWR.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4.5 l=0.35
**devattr s=26100,958 d=26100,958
R0 ctrl.n1 ctrl.t0 317.212
R1 ctrl.t0 ctrl.n0 317.212
R2 ctrl.n1 ctrl.t1 317.185
R3 ctrl.t1 ctrl.n0 317.185
R4 ctrl.n3 ctrl.t2 231.677
R5 ctrl.n2 ctrl.n1 68.35
R6 ctrl.n2 ctrl.n0 66.8028
R7 ctrl ctrl.n3 9.07858
R8 ctrl.n3 ctrl.n2 0.387869
R9 a_264_2813.n9 a_264_2813.t22 515.574
R10 a_264_2813.n4 a_264_2813.t22 515.574
R11 a_264_2813.n13 a_264_2813.n12 1.57443
R12 a_264_2813.t12 a_264_2813.n12 256.827
R13 a_264_2813.n13 a_264_2813.t21 515.226
R14 a_264_2813.t21 a_264_2813.n11 515.226
R15 a_264_2813.t3 a_264_2813.n1 515.226
R16 a_264_2813.n6 a_264_2813.t3 515.226
R17 a_264_2813.t6 a_264_2813.n1 515.226
R18 a_264_2813.n6 a_264_2813.t6 515.226
R19 a_264_2813.n1 a_264_2813.t17 515.226
R20 a_264_2813.t17 a_264_2813.n6 515.226
R21 a_264_2813.n1 a_264_2813.t18 515.226
R22 a_264_2813.t18 a_264_2813.n6 515.226
R23 a_264_2813.t26 a_264_2813.n0 515.226
R24 a_264_2813.n5 a_264_2813.t26 515.226
R25 a_264_2813.t5 a_264_2813.n0 515.226
R26 a_264_2813.n5 a_264_2813.t5 515.226
R27 a_264_2813.n0 a_264_2813.t16 515.226
R28 a_264_2813.t16 a_264_2813.n5 515.226
R29 a_264_2813.n0 a_264_2813.t24 515.226
R30 a_264_2813.t24 a_264_2813.n5 515.226
R31 a_264_2813.t25 a_264_2813.n2 515.226
R32 a_264_2813.n7 a_264_2813.t25 515.226
R33 a_264_2813.t4 a_264_2813.n2 515.226
R34 a_264_2813.n7 a_264_2813.t4 515.226
R35 a_264_2813.n2 a_264_2813.t15 515.226
R36 a_264_2813.t15 a_264_2813.n7 515.226
R37 a_264_2813.n2 a_264_2813.t8 515.226
R38 a_264_2813.t8 a_264_2813.n7 515.226
R39 a_264_2813.t9 a_264_2813.n3 515.226
R40 a_264_2813.n8 a_264_2813.t9 515.226
R41 a_264_2813.t13 a_264_2813.n3 515.226
R42 a_264_2813.n8 a_264_2813.t13 515.226
R43 a_264_2813.n3 a_264_2813.t23 515.226
R44 a_264_2813.t23 a_264_2813.n8 515.226
R45 a_264_2813.n3 a_264_2813.t7 515.226
R46 a_264_2813.t7 a_264_2813.n8 515.226
R47 a_264_2813.t10 a_264_2813.n4 515.226
R48 a_264_2813.n9 a_264_2813.t10 515.226
R49 a_264_2813.t19 a_264_2813.n4 515.226
R50 a_264_2813.n9 a_264_2813.t19 515.226
R51 a_264_2813.n17 a_264_2813.t14 317.212
R52 a_264_2813.t14 a_264_2813.n16 317.212
R53 a_264_2813.t20 a_264_2813.n16 317.185
R54 a_264_2813.n17 a_264_2813.t20 317.185
R55 a_264_2813.n10 a_264_2813.t11 231.684
R56 a_264_2813.n15 a_264_2813.n14 149.701
R57 a_264_2813.n10 a_264_2813.n16 68.09
R58 a_264_2813.n10 a_264_2813.n17 67.0628
R59 a_264_2813.t0 a_264_2813.n18 62.2152
R60 a_264_2813.n14 a_264_2813.t1 21.6705
R61 a_264_2813.n14 a_264_2813.t2 21.6705
R62 a_264_2813.n15 a_264_2813.n11 6.30606
R63 a_264_2813.n18 a_264_2813.n10 5.22455
R64 a_264_2813.n11 a_264_2813.n6 1.74235
R65 a_264_2813.n11 a_264_2813.n12 1.57443
R66 a_264_2813.n7 a_264_2813.n8 1.3918
R67 a_264_2813.n5 a_264_2813.n7 1.3918
R68 a_264_2813.n6 a_264_2813.n5 1.3918
R69 a_264_2813.n2 a_264_2813.n3 1.3918
R70 a_264_2813.n0 a_264_2813.n2 1.3918
R71 a_264_2813.n1 a_264_2813.n0 1.3918
R72 a_264_2813.n13 a_264_2813.n1 1.3918
R73 a_264_2813.n3 a_264_2813.n4 1.04398
R74 a_264_2813.n8 a_264_2813.n9 1.04398
R75 a_264_2813.n18 a_264_2813.n15 1.02596
R76 VPWR.n14 VPWR.n11 7260
R77 VPWR.n15 VPWR.n11 7260
R78 VPWR.n14 VPWR.n12 7260
R79 VPWR.n15 VPWR.n12 7260
R80 VPWR.n27 VPWR.n4 1796.47
R81 VPWR.n20 VPWR.n19 1796.47
R82 VPWR.n19 VPWR.n8 1796.47
R83 VPWR.n29 VPWR.n4 1796.47
R84 VPWR.n23 VPWR.n6 1055.29
R85 VPWR.n23 VPWR.n5 1055.29
R86 VPWR.n16 VPWR.n10 774.4
R87 VPWR.n13 VPWR.n10 774.4
R88 VPWR.n27 VPWR.n6 741.178
R89 VPWR.n20 VPWR.n6 741.178
R90 VPWR.n29 VPWR.n5 741.178
R91 VPWR.n8 VPWR.n5 741.178
R92 VPWR.t13 VPWR.n4 234.965
R93 VPWR.n19 VPWR.t25 234.965
R94 VPWR.n17 VPWR.n16 225.506
R95 VPWR.n13 VPWR.n0 225.506
R96 VPWR.n22 VPWR.t6 208.537
R97 VPWR.n22 VPWR.t27 208.537
R98 VPWR.n18 VPWR.n7 191.625
R99 VPWR.n26 VPWR.n2 191.625
R100 VPWR.n33 VPWR.t26 174.149
R101 VPWR.n33 VPWR.t28 174.053
R102 VPWR.n34 VPWR.t7 174.053
R103 VPWR.n35 VPWR.t14 174.053
R104 VPWR.t4 VPWR.n14 137.946
R105 VPWR.n15 VPWR.t16 137.946
R106 VPWR.n18 VPWR.n17 129.999
R107 VPWR.n31 VPWR.n2 112.566
R108 VPWR.n25 VPWR.n24 112.566
R109 VPWR.n24 VPWR.n3 112.566
R110 VPWR.t8 VPWR.t4 90.8824
R111 VPWR.t17 VPWR.t8 90.8824
R112 VPWR.t20 VPWR.t17 90.8824
R113 VPWR.t3 VPWR.t20 90.8824
R114 VPWR.t15 VPWR.t3 90.8824
R115 VPWR.t18 VPWR.t15 90.8824
R116 VPWR.t19 VPWR.t18 90.8824
R117 VPWR.t12 VPWR.t19 90.8824
R118 VPWR.t23 VPWR.t12 90.8824
R119 VPWR.t1 VPWR.t23 90.8824
R120 VPWR.t2 VPWR.t1 90.8824
R121 VPWR.t11 VPWR.t2 90.8824
R122 VPWR.t22 VPWR.t11 90.8824
R123 VPWR.t0 VPWR.t22 90.8824
R124 VPWR.t9 VPWR.t0 90.8824
R125 VPWR.t10 VPWR.t9 90.8824
R126 VPWR.t21 VPWR.t10 90.8824
R127 VPWR.t24 VPWR.t21 90.8824
R128 VPWR.t5 VPWR.t24 90.8824
R129 VPWR.t16 VPWR.t5 90.8824
R130 VPWR.n26 VPWR.n25 79.0593
R131 VPWR.n25 VPWR.n7 79.0593
R132 VPWR.n28 VPWR.t13 61.7891
R133 VPWR.n28 VPWR.t6 61.7891
R134 VPWR.t27 VPWR.n21 61.7891
R135 VPWR.n21 VPWR.t25 61.7891
R136 VPWR.n1 VPWR.n0 57.6005
R137 VPWR.n27 VPWR.n26 46.2505
R138 VPWR.n28 VPWR.n27 46.2505
R139 VPWR.n20 VPWR.n7 46.2505
R140 VPWR.n21 VPWR.n20 46.2505
R141 VPWR.n9 VPWR.n8 46.2505
R142 VPWR.n21 VPWR.n8 46.2505
R143 VPWR.n30 VPWR.n29 46.2505
R144 VPWR.n29 VPWR.n28 46.2505
R145 VPWR.n32 VPWR.n31 30.8117
R146 VPWR.n19 VPWR.n18 26.4291
R147 VPWR.n4 VPWR.n2 26.4291
R148 VPWR.n24 VPWR.n23 26.4291
R149 VPWR.n23 VPWR.n22 26.4291
R150 VPWR.n16 VPWR.n15 11.563
R151 VPWR.n14 VPWR.n13 11.563
R152 VPWR.n37 VPWR.n0 10.8709
R153 VPWR.n31 VPWR.n30 6.78838
R154 VPWR.n30 VPWR.n3 6.78838
R155 VPWR.n9 VPWR.n3 6.78838
R156 VPWR.n12 VPWR.n10 4.5127
R157 VPWR.t1 VPWR.n12 4.5127
R158 VPWR.n11 VPWR.n1 4.5127
R159 VPWR.t1 VPWR.n11 4.5127
R160 VPWR.n38 VPWR.n37 2.2055
R161 VPWR.n32 VPWR.n1 0.909142
R162 VPWR.n37 VPWR.n36 0.901542
R163 VPWR.n17 VPWR.n9 0.711611
R164 VPWR.n38 VPWR 0.4846
R165 VPWR.n36 VPWR.n35 0.46925
R166 VPWR VPWR.n38 0.368667
R167 VPWR.n34 VPWR.n33 0.122375
R168 VPWR.n36 VPWR.n32 0.106182
R169 VPWR.n35 VPWR.n34 0.097375
R170 bus.n10 bus.t1 53.5778
R171 bus.n18 bus.n17 47.2902
R172 bus.n20 bus.n14 47.0712
R173 bus.n19 bus.n15 47.0712
R174 bus.n18 bus.n16 47.0712
R175 bus.n10 bus.n9 47.0712
R176 bus.n11 bus.n8 47.0712
R177 bus.n12 bus.n7 47.0712
R178 bus.n13 bus.n6 47.0712
R179 bus.n23 bus.n22 47.0712
R180 bus.n23 bus.n21 47.0712
R181 bus.n1 bus.t26 20.5349
R182 bus.n4 bus.n3 16.6683
R183 bus.n1 bus.n0 16.5083
R184 bus.n4 bus.n2 16.5083
R185 bus.n17 bus.t5 6.34828
R186 bus.n17 bus.t3 6.34828
R187 bus.n14 bus.t17 6.34828
R188 bus.n14 bus.t20 6.34828
R189 bus.n15 bus.t13 6.34828
R190 bus.n15 bus.t2 6.34828
R191 bus.n16 bus.t0 6.34828
R192 bus.n16 bus.t18 6.34828
R193 bus.n9 bus.t19 6.34828
R194 bus.n9 bus.t4 6.34828
R195 bus.n8 bus.t10 6.34828
R196 bus.n8 bus.t16 6.34828
R197 bus.n7 bus.t6 6.34828
R198 bus.n7 bus.t12 6.34828
R199 bus.n6 bus.t9 6.34828
R200 bus.n6 bus.t15 6.34828
R201 bus.n22 bus.t11 6.34828
R202 bus.n22 bus.t14 6.34828
R203 bus.n21 bus.t8 6.34828
R204 bus.n21 bus.t7 6.34828
R205 bus.n3 bus.t25 3.86717
R206 bus.n3 bus.t24 3.86717
R207 bus.n0 bus.t22 3.86717
R208 bus.n0 bus.t21 3.86717
R209 bus.n2 bus.t23 3.86717
R210 bus.n2 bus.t27 3.86717
R211 bus.n26 bus.n25 0.6825
R212 bus.n13 bus.n12 0.1605
R213 bus.n12 bus.n11 0.1605
R214 bus.n11 bus.n10 0.1605
R215 bus.n19 bus.n18 0.1605
R216 bus.n20 bus.n19 0.1605
R217 bus.n24 bus.n13 0.142375
R218 bus.n25 bus.n24 0.1255
R219 bus.n5 bus.n1 0.121125
R220 bus.n24 bus.n20 0.088625
R221 bus bus.n26 0.0527222
R222 bus.n26 bus 0.0527222
R223 bus.n5 bus.n4 0.039875
R224 bus.n24 bus.n23 0.03175
R225 bus.n25 bus.n5 0.028625
R226 mod.n25 mod.t4 52.4447
R227 mod.n16 mod.n15 47.2312
R228 mod.n18 mod.n12 47.0712
R229 mod.n17 mod.n13 47.0712
R230 mod.n16 mod.n14 47.0712
R231 mod.n24 mod.n6 47.0712
R232 mod.n23 mod.n7 47.0712
R233 mod.n22 mod.n8 47.0712
R234 mod.n21 mod.n9 47.0712
R235 mod.n20 mod.n10 47.0712
R236 mod.n19 mod.n11 47.0712
R237 mod.n4 mod.t22 20.5349
R238 mod.n2 mod.n1 16.6895
R239 mod.n4 mod.n3 16.5083
R240 mod.n2 mod.n0 16.5083
R241 mod.n12 mod.t18 6.34828
R242 mod.n12 mod.t0 6.34828
R243 mod.n13 mod.t7 6.34828
R244 mod.n13 mod.t8 6.34828
R245 mod.n14 mod.t17 6.34828
R246 mod.n14 mod.t20 6.34828
R247 mod.n15 mod.t5 6.34828
R248 mod.n15 mod.t12 6.34828
R249 mod.n6 mod.t6 6.34828
R250 mod.n6 mod.t13 6.34828
R251 mod.n7 mod.t16 6.34828
R252 mod.n7 mod.t3 6.34828
R253 mod.n8 mod.t11 6.34828
R254 mod.n8 mod.t14 6.34828
R255 mod.n9 mod.t15 6.34828
R256 mod.n9 mod.t10 6.34828
R257 mod.n10 mod.t19 6.34828
R258 mod.n10 mod.t1 6.34828
R259 mod.n11 mod.t2 6.34828
R260 mod.n11 mod.t9 6.34828
R261 mod.n1 mod.t21 3.86717
R262 mod.n1 mod.t24 3.86717
R263 mod.n3 mod.t26 3.86717
R264 mod.n3 mod.t27 3.86717
R265 mod.n0 mod.t23 3.86717
R266 mod.n0 mod.t25 3.86717
R267 mod.n26 mod.n25 1.30798
R268 mod.n26 mod.n5 0.369625
R269 mod.n27 mod.n26 0.3415
R270 mod.n25 mod.n24 0.25425
R271 mod.n18 mod.n17 0.1605
R272 mod.n17 mod.n16 0.1605
R273 mod.n19 mod.n18 0.134562
R274 mod.n5 mod.n4 0.126125
R275 mod.n24 mod.n23 0.0805
R276 mod.n23 mod.n22 0.0805
R277 mod.n22 mod.n21 0.0805
R278 mod.n21 mod.n20 0.0805
R279 mod.n20 mod.n19 0.0805
R280 mod mod.n27 0.0527222
R281 mod.n27 mod 0.0527222
R282 mod.n5 mod.n2 0.034875
R283 VGND.n17 VGND.n7 81177.1
R284 VGND.n11 VGND.n8 6674.82
R285 VGND.n15 VGND.n8 6674.82
R286 VGND.n11 VGND.n9 6674.82
R287 VGND.n15 VGND.n9 6674.82
R288 VGND.n27 VGND.n5 2595.76
R289 VGND.n28 VGND.n5 2595.76
R290 VGND.n32 VGND.n3 2595.76
R291 VGND.n20 VGND.n4 1680.29
R292 VGND.n29 VGND.n4 1680.29
R293 VGND.n27 VGND.n20 915.471
R294 VGND.n20 VGND.n3 915.471
R295 VGND.n29 VGND.n28 915.471
R296 VGND.n30 VGND.n29 915.471
R297 VGND.t0 VGND.n18 681.569
R298 VGND.t0 VGND.n19 681.569
R299 VGND.n19 VGND.t9 681.569
R300 VGND.n18 VGND.n17 677.255
R301 VGND.n17 VGND.n16 653.227
R302 VGND.n32 VGND.n31 543.638
R303 VGND.n12 VGND.n10 433.695
R304 VGND.n14 VGND.n10 433.695
R305 VGND.n13 VGND.n12 433.695
R306 VGND.n14 VGND.n13 433.695
R307 VGND.t2 VGND.n7 388.878
R308 VGND.n16 VGND.t3 388.878
R309 VGND.n30 VGND.n2 292.5
R310 VGND.n28 VGND.n6 292.5
R311 VGND.n28 VGND.t0 292.5
R312 VGND.n27 VGND.n26 292.5
R313 VGND.t0 VGND.n27 292.5
R314 VGND.n3 VGND.n1 292.5
R315 VGND.t9 VGND.n3 292.5
R316 VGND.t5 VGND.t2 279.642
R317 VGND.t4 VGND.t5 279.642
R318 VGND.t6 VGND.t4 279.642
R319 VGND.t6 VGND.t7 279.642
R320 VGND.t7 VGND.t8 279.642
R321 VGND.t8 VGND.t3 279.642
R322 VGND.n31 VGND.n30 207.823
R323 VGND.n33 VGND.n2 168.66
R324 VGND.n21 VGND.n6 168.66
R325 VGND.n34 VGND.n33 110.314
R326 VGND.n24 VGND.n23 109.177
R327 VGND.n25 VGND.n24 108.424
R328 VGND.n22 VGND.n21 108.424
R329 VGND.n24 VGND.n4 83.5719
R330 VGND.n19 VGND.n4 83.5719
R331 VGND.n33 VGND.n32 83.5719
R332 VGND.n21 VGND.n5 83.5719
R333 VGND.n18 VGND.n5 83.5719
R334 VGND.n0 VGND.t1 64.0037
R335 VGND.n36 VGND.t10 62.2777
R336 VGND.n22 VGND.n0 61.835
R337 VGND.n31 VGND.t9 61.2599
R338 VGND.n23 VGND.n6 59.4829
R339 VGND.n23 VGND.n2 59.4829
R340 VGND.n13 VGND.n9 41.7862
R341 VGND.n9 VGND.t6 41.7862
R342 VGND.n10 VGND.n8 41.7862
R343 VGND.t6 VGND.n8 41.7862
R344 VGND.n15 VGND.n14 36.563
R345 VGND.n16 VGND.n15 36.563
R346 VGND.n12 VGND.n11 36.563
R347 VGND.n11 VGND.n7 36.563
R348 VGND.n26 VGND.n22 6.09207
R349 VGND.n26 VGND.n25 6.09207
R350 VGND.n25 VGND.n1 6.09207
R351 VGND.n34 VGND.n1 4.20291
R352 VGND.n37 VGND.n36 1.7055
R353 VGND.n35 VGND.n34 1.03383
R354 VGND.n37 VGND 0.829267
R355 VGND.n36 VGND.n35 0.5005
R356 VGND.n35 VGND.n0 0.2005
R357 VGND VGND.n37 0.024
C0 VPWR ctrl 1.07036f
C1 mod ctrl 0.052081f
C2 ctrl bus 0.007757f
C3 mod VPWR 1.79432f
C4 VPWR bus 1.99929f
C5 mod bus 23.4702f
C6 a_680_3582# ctrl 0.167494f
C7 VPWR a_680_3582# 1.08351f
C8 mod a_680_3582# 1.3552f
C9 a_680_3582# bus 0.687796f
.ends

