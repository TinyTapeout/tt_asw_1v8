magic
tech sky130A
magscale 1 2
timestamp 1711022820
<< error_p >>
rect -269 331 -211 337
rect -77 331 -19 337
rect 115 331 173 337
rect 307 331 365 337
rect -269 297 -257 331
rect -77 297 -65 331
rect 115 297 127 331
rect 307 297 319 331
rect -269 291 -211 297
rect -77 291 -19 297
rect 115 291 173 297
rect 307 291 365 297
rect -365 -297 -307 -291
rect -173 -297 -115 -291
rect 19 -297 77 -291
rect 211 -297 269 -291
rect -365 -331 -353 -297
rect -173 -331 -161 -297
rect 19 -331 31 -297
rect 211 -331 223 -297
rect -365 -337 -307 -331
rect -173 -337 -115 -331
rect 19 -337 77 -331
rect 211 -337 269 -331
<< nwell >>
rect -551 -469 551 469
<< pmos >>
rect -351 -250 -321 250
rect -255 -250 -225 250
rect -159 -250 -129 250
rect -63 -250 -33 250
rect 33 -250 63 250
rect 129 -250 159 250
rect 225 -250 255 250
rect 321 -250 351 250
<< pdiff >>
rect -413 238 -351 250
rect -413 -238 -401 238
rect -367 -238 -351 238
rect -413 -250 -351 -238
rect -321 238 -255 250
rect -321 -238 -305 238
rect -271 -238 -255 238
rect -321 -250 -255 -238
rect -225 238 -159 250
rect -225 -238 -209 238
rect -175 -238 -159 238
rect -225 -250 -159 -238
rect -129 238 -63 250
rect -129 -238 -113 238
rect -79 -238 -63 238
rect -129 -250 -63 -238
rect -33 238 33 250
rect -33 -238 -17 238
rect 17 -238 33 238
rect -33 -250 33 -238
rect 63 238 129 250
rect 63 -238 79 238
rect 113 -238 129 238
rect 63 -250 129 -238
rect 159 238 225 250
rect 159 -238 175 238
rect 209 -238 225 238
rect 159 -250 225 -238
rect 255 238 321 250
rect 255 -238 271 238
rect 305 -238 321 238
rect 255 -250 321 -238
rect 351 238 413 250
rect 351 -238 367 238
rect 401 -238 413 238
rect 351 -250 413 -238
<< pdiffc >>
rect -401 -238 -367 238
rect -305 -238 -271 238
rect -209 -238 -175 238
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
rect 175 -238 209 238
rect 271 -238 305 238
rect 367 -238 401 238
<< nsubdiff >>
rect -515 399 -419 433
rect 419 399 515 433
rect -515 337 -481 399
rect 481 337 515 399
rect -515 -399 -481 -337
rect 481 -399 515 -337
rect -515 -433 -419 -399
rect 419 -433 515 -399
<< nsubdiffcont >>
rect -419 399 419 433
rect -515 -337 -481 337
rect 481 -337 515 337
rect -419 -433 419 -399
<< poly >>
rect -273 331 -207 347
rect -273 297 -257 331
rect -223 297 -207 331
rect -273 281 -207 297
rect -81 331 -15 347
rect -81 297 -65 331
rect -31 297 -15 331
rect -81 281 -15 297
rect 111 331 177 347
rect 111 297 127 331
rect 161 297 177 331
rect 111 281 177 297
rect 303 331 369 347
rect 303 297 319 331
rect 353 297 369 331
rect 303 281 369 297
rect -351 250 -321 276
rect -255 250 -225 281
rect -159 250 -129 276
rect -63 250 -33 281
rect 33 250 63 276
rect 129 250 159 281
rect 225 250 255 276
rect 321 250 351 281
rect -351 -281 -321 -250
rect -255 -276 -225 -250
rect -159 -281 -129 -250
rect -63 -276 -33 -250
rect 33 -281 63 -250
rect 129 -276 159 -250
rect 225 -281 255 -250
rect 321 -276 351 -250
rect -369 -297 -303 -281
rect -369 -331 -353 -297
rect -319 -331 -303 -297
rect -369 -347 -303 -331
rect -177 -297 -111 -281
rect -177 -331 -161 -297
rect -127 -331 -111 -297
rect -177 -347 -111 -331
rect 15 -297 81 -281
rect 15 -331 31 -297
rect 65 -331 81 -297
rect 15 -347 81 -331
rect 207 -297 273 -281
rect 207 -331 223 -297
rect 257 -331 273 -297
rect 207 -347 273 -331
<< polycont >>
rect -257 297 -223 331
rect -65 297 -31 331
rect 127 297 161 331
rect 319 297 353 331
rect -353 -331 -319 -297
rect -161 -331 -127 -297
rect 31 -331 65 -297
rect 223 -331 257 -297
<< locali >>
rect -515 399 -419 433
rect 419 399 515 433
rect -515 337 -481 399
rect 481 337 515 399
rect -273 297 -257 331
rect -223 297 -207 331
rect -81 297 -65 331
rect -31 297 -15 331
rect 111 297 127 331
rect 161 297 177 331
rect 303 297 319 331
rect 353 297 369 331
rect -401 238 -367 254
rect -401 -254 -367 -238
rect -305 238 -271 254
rect -305 -254 -271 -238
rect -209 238 -175 254
rect -209 -254 -175 -238
rect -113 238 -79 254
rect -113 -254 -79 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 79 238 113 254
rect 79 -254 113 -238
rect 175 238 209 254
rect 175 -254 209 -238
rect 271 238 305 254
rect 271 -254 305 -238
rect 367 238 401 254
rect 367 -254 401 -238
rect -369 -331 -353 -297
rect -319 -331 -303 -297
rect -177 -331 -161 -297
rect -127 -331 -111 -297
rect 15 -331 31 -297
rect 65 -331 81 -297
rect 207 -331 223 -297
rect 257 -331 273 -297
rect -515 -399 -481 -337
rect 481 -399 515 -337
rect -515 -433 -419 -399
rect 419 -433 515 -399
<< viali >>
rect -257 297 -223 331
rect -65 297 -31 331
rect 127 297 161 331
rect 319 297 353 331
rect -401 -238 -367 238
rect -305 -238 -271 238
rect -209 -238 -175 238
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
rect 175 -238 209 238
rect 271 -238 305 238
rect 367 -238 401 238
rect -353 -331 -319 -297
rect -161 -331 -127 -297
rect 31 -331 65 -297
rect 223 -331 257 -297
<< metal1 >>
rect -269 331 -211 337
rect -269 297 -257 331
rect -223 297 -211 331
rect -269 291 -211 297
rect -77 331 -19 337
rect -77 297 -65 331
rect -31 297 -19 331
rect -77 291 -19 297
rect 115 331 173 337
rect 115 297 127 331
rect 161 297 173 331
rect 115 291 173 297
rect 307 331 365 337
rect 307 297 319 331
rect 353 297 365 331
rect 307 291 365 297
rect -407 238 -361 250
rect -407 -238 -401 238
rect -367 -238 -361 238
rect -407 -250 -361 -238
rect -311 238 -265 250
rect -311 -238 -305 238
rect -271 -238 -265 238
rect -311 -250 -265 -238
rect -215 238 -169 250
rect -215 -238 -209 238
rect -175 -238 -169 238
rect -215 -250 -169 -238
rect -119 238 -73 250
rect -119 -238 -113 238
rect -79 -238 -73 238
rect -119 -250 -73 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 73 238 119 250
rect 73 -238 79 238
rect 113 -238 119 238
rect 73 -250 119 -238
rect 169 238 215 250
rect 169 -238 175 238
rect 209 -238 215 238
rect 169 -250 215 -238
rect 265 238 311 250
rect 265 -238 271 238
rect 305 -238 311 238
rect 265 -250 311 -238
rect 361 238 407 250
rect 361 -238 367 238
rect 401 -238 407 238
rect 361 -250 407 -238
rect -365 -297 -307 -291
rect -365 -331 -353 -297
rect -319 -331 -307 -297
rect -365 -337 -307 -331
rect -173 -297 -115 -291
rect -173 -331 -161 -297
rect -127 -331 -115 -297
rect -173 -337 -115 -331
rect 19 -297 77 -291
rect 19 -331 31 -297
rect 65 -331 77 -297
rect 19 -337 77 -331
rect 211 -297 269 -291
rect 211 -331 223 -297
rect 257 -331 269 -297
rect 211 -337 269 -331
<< properties >>
string FIXED_BBOX -498 -416 498 416
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
