magic
tech sky130A
magscale 1 2
timestamp 1711022820
<< error_p >>
rect -77 322 -19 328
rect 115 322 173 328
rect -77 288 -65 322
rect 115 288 127 322
rect -77 282 -19 288
rect 115 282 173 288
rect -173 -288 -115 -282
rect 19 -288 77 -282
rect -173 -322 -161 -288
rect 19 -322 31 -288
rect -173 -328 -115 -322
rect 19 -328 77 -322
<< pwell >>
rect -359 -460 359 460
<< nmos >>
rect -159 -250 -129 250
rect -63 -250 -33 250
rect 33 -250 63 250
rect 129 -250 159 250
<< ndiff >>
rect -221 238 -159 250
rect -221 -238 -209 238
rect -175 -238 -159 238
rect -221 -250 -159 -238
rect -129 238 -63 250
rect -129 -238 -113 238
rect -79 -238 -63 238
rect -129 -250 -63 -238
rect -33 238 33 250
rect -33 -238 -17 238
rect 17 -238 33 238
rect -33 -250 33 -238
rect 63 238 129 250
rect 63 -238 79 238
rect 113 -238 129 238
rect 63 -250 129 -238
rect 159 238 221 250
rect 159 -238 175 238
rect 209 -238 221 238
rect 159 -250 221 -238
<< ndiffc >>
rect -209 -238 -175 238
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
rect 175 -238 209 238
<< psubdiff >>
rect -323 390 -227 424
rect 227 390 323 424
rect -323 328 -289 390
rect 289 328 323 390
rect -323 -390 -289 -328
rect 289 -390 323 -328
rect -323 -424 -227 -390
rect 227 -424 323 -390
<< psubdiffcont >>
rect -227 390 227 424
rect -323 -328 -289 328
rect 289 -328 323 328
rect -227 -424 227 -390
<< poly >>
rect -81 322 -15 338
rect -81 288 -65 322
rect -31 288 -15 322
rect -159 250 -129 276
rect -81 272 -15 288
rect 111 322 177 338
rect 111 288 127 322
rect 161 288 177 322
rect -63 250 -33 272
rect 33 250 63 276
rect 111 272 177 288
rect 129 250 159 272
rect -159 -272 -129 -250
rect -177 -288 -111 -272
rect -63 -276 -33 -250
rect 33 -272 63 -250
rect -177 -322 -161 -288
rect -127 -322 -111 -288
rect -177 -338 -111 -322
rect 15 -288 81 -272
rect 129 -276 159 -250
rect 15 -322 31 -288
rect 65 -322 81 -288
rect 15 -338 81 -322
<< polycont >>
rect -65 288 -31 322
rect 127 288 161 322
rect -161 -322 -127 -288
rect 31 -322 65 -288
<< locali >>
rect -323 390 -227 424
rect 227 390 323 424
rect -323 328 -289 390
rect 289 328 323 390
rect -81 288 -65 322
rect -31 288 -15 322
rect 111 288 127 322
rect 161 288 177 322
rect -209 238 -175 254
rect -209 -254 -175 -238
rect -113 238 -79 254
rect -113 -254 -79 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 79 238 113 254
rect 79 -254 113 -238
rect 175 238 209 254
rect 175 -254 209 -238
rect -177 -322 -161 -288
rect -127 -322 -111 -288
rect 15 -322 31 -288
rect 65 -322 81 -288
rect -323 -390 -289 -328
rect 289 -390 323 -328
rect -323 -424 -227 -390
rect 227 -424 323 -390
<< viali >>
rect -65 288 -31 322
rect 127 288 161 322
rect -209 -238 -175 238
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
rect 175 -238 209 238
rect -161 -322 -127 -288
rect 31 -322 65 -288
<< metal1 >>
rect -77 322 -19 328
rect -77 288 -65 322
rect -31 288 -19 322
rect -77 282 -19 288
rect 115 322 173 328
rect 115 288 127 322
rect 161 288 173 322
rect 115 282 173 288
rect -215 238 -169 250
rect -215 -238 -209 238
rect -175 -238 -169 238
rect -215 -250 -169 -238
rect -119 238 -73 250
rect -119 -238 -113 238
rect -79 -238 -73 238
rect -119 -250 -73 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 73 238 119 250
rect 73 -238 79 238
rect 113 -238 119 238
rect 73 -250 119 -238
rect 169 238 215 250
rect 169 -238 175 238
rect 209 -238 215 238
rect 169 -250 215 -238
rect -173 -288 -115 -282
rect -173 -322 -161 -288
rect -127 -322 -115 -288
rect -173 -328 -115 -322
rect 19 -288 77 -282
rect 19 -322 31 -288
rect 65 -322 77 -288
rect 19 -328 77 -322
<< properties >>
string FIXED_BBOX -306 -407 306 407
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
