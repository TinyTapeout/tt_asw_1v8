** sch_path: /home/matt/work/asic-workshop/shuttle-2404/tt-analog-switch/xschem/tt_asw_1v8.sch
.subckt tt_asw_1v8 VPWR ctrl mod bus VGND
*.PININFO VPWR:B VGND:B mod:B bus:B ctrl:I
XM4 tgon tgon_n VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 m=1
XM3 tgon tgon_n VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=2 m=1
XM2 tgon_n ctrl VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 m=1
XM1 tgon_n ctrl VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=2 m=1
XM6 bus tgon mod VGND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=12 nf=4 m=1
XM5 bus tgon_n mod VPWR sky130_fd_pr__pfet_01v8_lvt L=0.5 W=21 nf=7 m=1
.ends
.end
