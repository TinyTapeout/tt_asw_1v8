magic
tech sky130A
magscale 1 2
timestamp 1712309281
<< pwell >>
rect -483 -510 483 510
<< nmoslvt >>
rect -287 -300 -187 300
rect -129 -300 -29 300
rect 29 -300 129 300
rect 187 -300 287 300
<< ndiff >>
rect -345 288 -287 300
rect -345 -288 -333 288
rect -299 -288 -287 288
rect -345 -300 -287 -288
rect -187 288 -129 300
rect -187 -288 -175 288
rect -141 -288 -129 288
rect -187 -300 -129 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 129 288 187 300
rect 129 -288 141 288
rect 175 -288 187 288
rect 129 -300 187 -288
rect 287 288 345 300
rect 287 -288 299 288
rect 333 -288 345 288
rect 287 -300 345 -288
<< ndiffc >>
rect -333 -288 -299 288
rect -175 -288 -141 288
rect -17 -288 17 288
rect 141 -288 175 288
rect 299 -288 333 288
<< psubdiff >>
rect -447 440 -351 474
rect 351 440 447 474
rect -447 378 -413 440
rect 413 378 447 440
rect -447 -440 -413 -378
rect 413 -440 447 -378
rect -447 -474 -351 -440
rect 351 -474 447 -440
<< psubdiffcont >>
rect -351 440 351 474
rect -447 -378 -413 378
rect 413 -378 447 378
rect -351 -474 351 -440
<< poly >>
rect -287 372 -187 388
rect -287 338 -271 372
rect -203 338 -187 372
rect -287 300 -187 338
rect -129 372 -29 388
rect -129 338 -113 372
rect -45 338 -29 372
rect -129 300 -29 338
rect 29 372 129 388
rect 29 338 45 372
rect 113 338 129 372
rect 29 300 129 338
rect 187 372 287 388
rect 187 338 203 372
rect 271 338 287 372
rect 187 300 287 338
rect -287 -338 -187 -300
rect -287 -372 -271 -338
rect -203 -372 -187 -338
rect -287 -388 -187 -372
rect -129 -338 -29 -300
rect -129 -372 -113 -338
rect -45 -372 -29 -338
rect -129 -388 -29 -372
rect 29 -338 129 -300
rect 29 -372 45 -338
rect 113 -372 129 -338
rect 29 -388 129 -372
rect 187 -338 287 -300
rect 187 -372 203 -338
rect 271 -372 287 -338
rect 187 -388 287 -372
<< polycont >>
rect -271 338 -203 372
rect -113 338 -45 372
rect 45 338 113 372
rect 203 338 271 372
rect -271 -372 -203 -338
rect -113 -372 -45 -338
rect 45 -372 113 -338
rect 203 -372 271 -338
<< locali >>
rect -447 440 -351 474
rect 351 440 447 474
rect -447 378 -413 440
rect 413 378 447 440
rect -287 338 -271 372
rect -203 338 -187 372
rect -129 338 -113 372
rect -45 338 -29 372
rect 29 338 45 372
rect 113 338 129 372
rect 187 338 203 372
rect 271 338 287 372
rect -333 288 -299 304
rect -333 -304 -299 -288
rect -175 288 -141 304
rect -175 -304 -141 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 141 288 175 304
rect 141 -304 175 -288
rect 299 288 333 304
rect 299 -304 333 -288
rect -287 -372 -271 -338
rect -203 -372 -187 -338
rect -129 -372 -113 -338
rect -45 -372 -29 -338
rect 29 -372 45 -338
rect 113 -372 129 -338
rect 187 -372 203 -338
rect 271 -372 287 -338
rect -447 -440 -413 -378
rect 413 -440 447 -378
rect -447 -474 -351 -440
rect 351 -474 447 -440
<< viali >>
rect -271 338 -203 372
rect -113 338 -45 372
rect 45 338 113 372
rect 203 338 271 372
rect -333 -288 -299 288
rect -175 -288 -141 288
rect -17 -288 17 288
rect 141 -288 175 288
rect 299 -288 333 288
rect -271 -372 -203 -338
rect -113 -372 -45 -338
rect 45 -372 113 -338
rect 203 -372 271 -338
<< metal1 >>
rect -283 372 -191 378
rect -283 338 -271 372
rect -203 338 -191 372
rect -283 332 -191 338
rect -125 372 -33 378
rect -125 338 -113 372
rect -45 338 -33 372
rect -125 332 -33 338
rect 33 372 125 378
rect 33 338 45 372
rect 113 338 125 372
rect 33 332 125 338
rect 191 372 283 378
rect 191 338 203 372
rect 271 338 283 372
rect 191 332 283 338
rect -339 288 -293 300
rect -339 -288 -333 288
rect -299 -288 -293 288
rect -339 -300 -293 -288
rect -181 288 -135 300
rect -181 -288 -175 288
rect -141 -288 -135 288
rect -181 -300 -135 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 135 288 181 300
rect 135 -288 141 288
rect 175 -288 181 288
rect 135 -300 181 -288
rect 293 288 339 300
rect 293 -288 299 288
rect 333 -288 339 288
rect 293 -300 339 -288
rect -283 -338 -191 -332
rect -283 -372 -271 -338
rect -203 -372 -191 -338
rect -283 -378 -191 -372
rect -125 -338 -33 -332
rect -125 -372 -113 -338
rect -45 -372 -33 -338
rect -125 -378 -33 -372
rect 33 -338 125 -332
rect 33 -372 45 -338
rect 113 -372 125 -338
rect 33 -378 125 -372
rect 191 -338 283 -332
rect 191 -372 203 -338
rect 271 -372 283 -338
rect 191 -378 283 -372
<< properties >>
string FIXED_BBOX -430 -457 430 457
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 3 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
