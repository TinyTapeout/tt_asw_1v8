VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_asw_1v8
  CLASS BLOCK ;
  FOREIGN tt_asw_1v8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.400 BY 21.760 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.600 0.000 1.800 21.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.600 0.000 17.800 21.760 ;
    END
  END VPWR
  PIN mod
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 6.090000 ;
    PORT
      LAYER met4 ;
        RECT 8.750 19.760 9.650 21.760 ;
    END
  END mod
  PIN bus
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 5.220000 ;
    PORT
      LAYER met4 ;
        RECT 8.750 11.760 9.650 13.760 ;
    END
  END bus
  PIN ctrl
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met3 ;
        RECT 4.450 20.860 4.750 21.760 ;
    END
  END ctrl
  OBS
      LAYER pwell ;
        RECT 0.690 16.860 4.380 20.460 ;
      LAYER nwell ;
        RECT 0.170 12.970 4.900 16.660 ;
      LAYER pwell ;
        RECT 4.900 14.200 9.730 19.300 ;
      LAYER nwell ;
        RECT 9.800 14.150 17.000 19.340 ;
      LAYER li1 ;
        RECT 0.600 20.100 17.800 21.760 ;
        RECT 0.870 17.210 1.040 20.100 ;
        RECT 1.580 19.600 1.910 19.770 ;
        RECT 1.440 17.890 1.610 19.430 ;
        RECT 1.880 17.890 2.050 19.430 ;
        RECT 1.580 17.550 1.910 17.720 ;
        RECT 2.450 17.210 2.620 20.100 ;
        RECT 3.160 19.600 3.490 19.770 ;
        RECT 3.020 17.890 3.190 19.430 ;
        RECT 3.460 17.890 3.630 19.430 ;
        RECT 3.160 17.550 3.490 17.720 ;
        RECT 4.030 17.210 4.200 20.100 ;
        RECT 0.870 17.040 4.200 17.210 ;
        RECT 5.080 18.950 9.550 20.100 ;
        RECT 0.350 16.310 4.720 16.480 ;
        RECT 0.350 13.320 0.520 16.310 ;
        RECT 1.075 15.795 1.895 15.975 ;
        RECT 0.920 14.045 1.090 15.585 ;
        RECT 1.400 14.045 1.570 15.585 ;
        RECT 1.880 14.045 2.050 15.585 ;
        RECT 1.075 13.655 1.895 13.835 ;
        RECT 2.450 13.320 2.620 16.310 ;
        RECT 3.175 15.795 3.995 15.975 ;
        RECT 3.020 14.045 3.190 15.585 ;
        RECT 3.500 14.045 3.670 15.585 ;
        RECT 3.980 14.045 4.150 15.585 ;
        RECT 3.175 13.655 3.995 13.835 ;
        RECT 4.550 13.320 4.720 16.310 ;
        RECT 5.080 14.550 5.250 18.950 ;
        RECT 5.880 18.440 6.380 18.610 ;
        RECT 6.670 18.440 7.170 18.610 ;
        RECT 7.460 18.440 7.960 18.610 ;
        RECT 8.250 18.440 8.750 18.610 ;
        RECT 5.650 15.230 5.820 18.270 ;
        RECT 6.440 15.230 6.610 18.270 ;
        RECT 7.230 15.230 7.400 18.270 ;
        RECT 8.020 15.230 8.190 18.270 ;
        RECT 8.810 15.230 8.980 18.270 ;
        RECT 5.880 14.890 6.380 15.060 ;
        RECT 6.670 14.890 7.170 15.060 ;
        RECT 7.460 14.890 7.960 15.060 ;
        RECT 8.250 14.890 8.750 15.060 ;
        RECT 9.380 14.550 9.550 18.950 ;
        RECT 5.080 14.380 9.550 14.550 ;
        RECT 9.980 18.990 16.820 19.160 ;
        RECT 9.980 14.500 10.150 18.990 ;
        RECT 10.780 18.480 11.280 18.650 ;
        RECT 11.570 18.480 12.070 18.650 ;
        RECT 12.360 18.480 12.860 18.650 ;
        RECT 13.150 18.480 13.650 18.650 ;
        RECT 13.940 18.480 14.440 18.650 ;
        RECT 14.730 18.480 15.230 18.650 ;
        RECT 15.520 18.480 16.020 18.650 ;
        RECT 10.550 15.225 10.720 18.265 ;
        RECT 11.340 15.225 11.510 18.265 ;
        RECT 12.130 15.225 12.300 18.265 ;
        RECT 12.920 15.225 13.090 18.265 ;
        RECT 13.710 15.225 13.880 18.265 ;
        RECT 14.500 15.225 14.670 18.265 ;
        RECT 15.290 15.225 15.460 18.265 ;
        RECT 16.080 15.225 16.250 18.265 ;
        RECT 10.780 14.840 11.280 15.010 ;
        RECT 11.570 14.840 12.070 15.010 ;
        RECT 12.360 14.840 12.860 15.010 ;
        RECT 13.150 14.840 13.650 15.010 ;
        RECT 13.940 14.840 14.440 15.010 ;
        RECT 14.730 14.840 15.230 15.010 ;
        RECT 15.520 14.840 16.020 15.010 ;
        RECT 16.650 14.500 16.820 18.990 ;
        RECT 9.980 13.320 16.820 14.500 ;
        RECT 0.350 13.150 17.800 13.320 ;
        RECT 0.600 11.760 17.800 13.150 ;
      LAYER mcon ;
        RECT 0.700 20.660 1.700 21.660 ;
        RECT 2.000 20.610 17.700 20.780 ;
        RECT 1.660 19.600 1.830 19.770 ;
        RECT 1.440 17.970 1.610 19.350 ;
        RECT 1.880 17.970 2.050 19.350 ;
        RECT 1.660 17.550 1.830 17.720 ;
        RECT 3.240 19.600 3.410 19.770 ;
        RECT 3.020 17.970 3.190 19.350 ;
        RECT 3.460 17.970 3.630 19.350 ;
        RECT 3.240 17.550 3.410 17.720 ;
        RECT 1.160 15.800 1.330 15.970 ;
        RECT 1.640 15.800 1.810 15.970 ;
        RECT 0.920 14.125 1.090 15.505 ;
        RECT 1.400 14.125 1.570 15.505 ;
        RECT 1.880 14.125 2.050 15.505 ;
        RECT 1.160 13.660 1.330 13.830 ;
        RECT 1.640 13.660 1.810 13.830 ;
        RECT 3.260 15.800 3.430 15.970 ;
        RECT 3.740 15.800 3.910 15.970 ;
        RECT 3.020 14.125 3.190 15.505 ;
        RECT 3.500 14.125 3.670 15.505 ;
        RECT 3.980 14.125 4.150 15.505 ;
        RECT 3.260 13.660 3.430 13.830 ;
        RECT 3.740 13.660 3.910 13.830 ;
        RECT 5.960 18.440 6.300 18.610 ;
        RECT 6.750 18.440 7.090 18.610 ;
        RECT 7.540 18.440 7.880 18.610 ;
        RECT 8.330 18.440 8.670 18.610 ;
        RECT 5.650 15.310 5.820 18.190 ;
        RECT 6.440 15.310 6.610 18.190 ;
        RECT 7.230 15.310 7.400 18.190 ;
        RECT 8.020 15.310 8.190 18.190 ;
        RECT 8.810 15.310 8.980 18.190 ;
        RECT 5.960 14.890 6.300 15.060 ;
        RECT 6.750 14.890 7.090 15.060 ;
        RECT 7.540 14.890 7.880 15.060 ;
        RECT 8.330 14.890 8.670 15.060 ;
        RECT 10.860 18.480 11.200 18.650 ;
        RECT 11.650 18.480 11.990 18.650 ;
        RECT 12.440 18.480 12.780 18.650 ;
        RECT 13.230 18.480 13.570 18.650 ;
        RECT 14.020 18.480 14.360 18.650 ;
        RECT 14.810 18.480 15.150 18.650 ;
        RECT 15.600 18.480 15.940 18.650 ;
        RECT 10.550 15.305 10.720 18.185 ;
        RECT 11.340 15.305 11.510 18.185 ;
        RECT 12.130 15.305 12.300 18.185 ;
        RECT 12.920 15.305 13.090 18.185 ;
        RECT 13.710 15.305 13.880 18.185 ;
        RECT 14.500 15.305 14.670 18.185 ;
        RECT 15.290 15.305 15.460 18.185 ;
        RECT 16.080 15.305 16.250 18.185 ;
        RECT 10.860 14.840 11.200 15.010 ;
        RECT 11.650 14.840 11.990 15.010 ;
        RECT 12.440 14.840 12.780 15.010 ;
        RECT 13.230 14.840 13.570 15.010 ;
        RECT 14.020 14.840 14.360 15.010 ;
        RECT 14.810 14.840 15.150 15.010 ;
        RECT 15.600 14.840 15.940 15.010 ;
        RECT 0.700 12.740 16.400 12.910 ;
        RECT 16.700 11.860 17.700 12.860 ;
      LAYER met1 ;
        RECT 0.600 20.560 17.800 21.760 ;
        RECT 0.950 19.560 1.890 19.810 ;
        RECT 2.530 19.560 3.470 19.810 ;
        RECT 0.950 17.760 1.180 19.560 ;
        RECT 1.410 17.910 1.670 19.410 ;
        RECT 1.820 17.910 2.080 19.410 ;
        RECT 2.530 17.760 2.760 19.560 ;
        RECT 2.990 17.910 3.250 19.410 ;
        RECT 3.400 17.910 3.660 19.410 ;
        RECT 5.140 18.410 8.730 18.640 ;
        RECT 10.040 18.450 16.020 18.680 ;
        RECT 0.950 17.510 1.890 17.760 ;
        RECT 2.530 17.510 3.470 17.760 ;
        RECT 0.950 16.940 1.180 17.510 ;
        RECT 0.920 16.580 1.210 16.940 ;
        RECT 2.530 16.920 2.760 17.510 ;
        RECT 5.140 16.920 5.370 18.410 ;
        RECT 2.510 16.860 2.780 16.920 ;
        RECT 2.510 16.660 4.700 16.860 ;
        RECT 2.510 16.600 2.780 16.660 ;
        RECT 0.950 16.010 1.180 16.580 ;
        RECT 2.530 16.010 2.760 16.600 ;
        RECT 0.430 15.760 1.900 16.010 ;
        RECT 2.530 15.760 4.000 16.010 ;
        RECT 0.430 13.870 0.660 15.760 ;
        RECT 0.890 14.060 1.150 15.570 ;
        RECT 1.350 14.060 1.620 15.570 ;
        RECT 1.820 14.060 2.080 15.570 ;
        RECT 2.530 13.870 2.760 15.760 ;
        RECT 2.990 14.060 3.250 15.570 ;
        RECT 3.450 14.060 3.720 15.570 ;
        RECT 3.920 14.060 4.180 15.570 ;
        RECT 4.500 14.600 4.700 16.660 ;
        RECT 5.120 16.600 5.390 16.920 ;
        RECT 5.140 15.090 5.370 16.600 ;
        RECT 5.600 15.240 5.870 18.250 ;
        RECT 6.390 15.240 6.660 18.250 ;
        RECT 7.180 15.240 7.450 18.250 ;
        RECT 7.970 15.240 8.240 18.250 ;
        RECT 8.760 15.240 9.030 18.250 ;
        RECT 10.040 16.860 10.270 18.450 ;
        RECT 9.500 16.660 10.270 16.860 ;
        RECT 5.140 14.860 8.730 15.090 ;
        RECT 9.500 14.600 9.700 16.660 ;
        RECT 10.040 15.040 10.270 16.660 ;
        RECT 10.500 15.240 10.770 18.250 ;
        RECT 11.290 15.240 11.560 18.250 ;
        RECT 12.080 15.240 12.350 18.250 ;
        RECT 12.870 15.240 13.140 18.250 ;
        RECT 13.660 15.240 13.930 18.250 ;
        RECT 14.450 15.240 14.720 18.250 ;
        RECT 15.240 15.240 15.510 18.250 ;
        RECT 16.030 15.240 16.300 18.250 ;
        RECT 10.040 14.810 16.020 15.040 ;
        RECT 4.500 14.400 9.700 14.600 ;
        RECT 0.430 13.620 1.900 13.870 ;
        RECT 2.530 13.620 4.000 13.870 ;
        RECT 0.600 11.760 17.800 12.960 ;
      LAYER via ;
        RECT 0.700 20.660 1.700 21.660 ;
        RECT 2.990 20.660 3.250 21.660 ;
        RECT 1.410 17.940 1.670 19.380 ;
        RECT 1.820 17.940 2.080 19.380 ;
        RECT 2.990 17.940 3.250 19.380 ;
        RECT 3.400 17.940 3.660 19.380 ;
        RECT 0.920 16.610 1.210 16.910 ;
        RECT 2.510 16.630 2.780 16.890 ;
        RECT 0.890 14.090 1.150 15.540 ;
        RECT 1.350 14.090 1.620 15.540 ;
        RECT 1.820 14.090 2.080 15.540 ;
        RECT 2.990 14.090 3.250 15.540 ;
        RECT 3.450 14.090 3.720 15.540 ;
        RECT 3.920 14.090 4.180 15.540 ;
        RECT 5.120 16.630 5.390 16.890 ;
        RECT 5.600 15.280 5.870 18.210 ;
        RECT 6.390 15.280 6.660 18.210 ;
        RECT 7.180 15.280 7.450 18.210 ;
        RECT 7.970 15.280 8.240 18.210 ;
        RECT 8.760 15.280 9.030 18.210 ;
        RECT 10.500 15.280 10.770 18.210 ;
        RECT 11.290 15.280 11.560 18.210 ;
        RECT 12.080 15.280 12.350 18.210 ;
        RECT 12.870 15.280 13.140 18.210 ;
        RECT 13.660 15.280 13.930 18.210 ;
        RECT 14.450 15.280 14.720 18.210 ;
        RECT 15.240 15.280 15.510 18.210 ;
        RECT 16.030 15.280 16.300 18.210 ;
        RECT 0.890 11.860 1.150 12.860 ;
        RECT 1.820 11.860 2.080 12.860 ;
        RECT 2.990 11.860 3.250 12.860 ;
        RECT 3.920 11.860 4.180 12.860 ;
        RECT 16.700 11.860 17.700 12.860 ;
      LAYER met2 ;
        RECT 0.600 20.560 1.800 21.760 ;
        RECT 1.410 17.910 1.670 20.560 ;
        RECT 0.920 16.560 1.210 16.960 ;
        RECT 1.820 16.860 2.080 19.410 ;
        RECT 2.990 17.910 3.250 21.760 ;
        RECT 2.480 16.860 2.810 16.890 ;
        RECT 1.350 16.660 2.810 16.860 ;
        RECT 3.400 16.860 3.660 19.410 ;
        RECT 5.090 16.860 5.420 16.890 ;
        RECT 3.400 16.660 5.420 16.860 ;
        RECT 0.890 11.760 1.150 15.570 ;
        RECT 1.350 14.060 1.620 16.660 ;
        RECT 2.480 16.630 2.810 16.660 ;
        RECT 1.820 11.760 2.080 15.570 ;
        RECT 2.990 11.760 3.250 15.570 ;
        RECT 3.450 14.060 3.720 16.660 ;
        RECT 5.090 16.630 5.420 16.660 ;
        RECT 3.920 11.760 4.180 15.570 ;
        RECT 5.590 15.230 5.880 18.260 ;
        RECT 6.380 15.230 6.670 18.260 ;
        RECT 7.170 15.230 7.460 18.260 ;
        RECT 7.960 15.230 8.250 18.260 ;
        RECT 8.750 15.230 9.040 18.260 ;
        RECT 10.490 15.230 10.780 18.260 ;
        RECT 11.280 15.230 11.570 18.260 ;
        RECT 12.070 15.230 12.360 18.260 ;
        RECT 12.860 15.230 13.150 18.260 ;
        RECT 13.650 15.230 13.940 18.260 ;
        RECT 14.440 15.230 14.730 18.260 ;
        RECT 15.230 15.230 15.520 18.260 ;
        RECT 16.020 15.230 16.310 18.260 ;
        RECT 16.600 11.760 17.800 12.960 ;
      LAYER via2 ;
        RECT 0.700 20.660 1.700 21.660 ;
        RECT 0.920 16.610 1.210 16.910 ;
        RECT 5.590 15.280 5.880 18.210 ;
        RECT 6.380 15.280 6.670 18.210 ;
        RECT 7.170 15.280 7.460 18.210 ;
        RECT 7.960 15.280 8.250 18.210 ;
        RECT 8.750 15.280 9.040 18.210 ;
        RECT 10.490 15.280 10.780 18.210 ;
        RECT 11.280 15.280 11.570 18.210 ;
        RECT 12.070 15.280 12.360 18.210 ;
        RECT 12.860 15.280 13.150 18.210 ;
        RECT 13.650 15.280 13.940 18.210 ;
        RECT 14.440 15.280 14.730 18.210 ;
        RECT 15.230 15.280 15.520 18.210 ;
        RECT 16.020 15.280 16.310 18.210 ;
        RECT 16.700 11.860 17.700 12.860 ;
      LAYER met3 ;
        RECT 0.600 20.560 1.800 21.760 ;
        RECT 0.890 16.910 1.240 16.940 ;
        RECT 4.450 16.910 4.750 20.860 ;
        RECT 8.750 19.760 9.650 21.760 ;
        RECT 0.890 16.610 4.750 16.910 ;
        RECT 5.560 18.700 15.550 19.760 ;
        RECT 0.890 16.580 1.240 16.610 ;
        RECT 5.560 15.250 5.910 18.700 ;
        RECT 6.350 14.790 6.700 18.240 ;
        RECT 7.140 15.250 7.490 18.700 ;
        RECT 7.930 14.790 8.280 18.240 ;
        RECT 8.720 15.250 9.070 18.700 ;
        RECT 10.460 15.250 10.810 18.700 ;
        RECT 11.250 14.790 11.600 18.240 ;
        RECT 12.040 15.250 12.390 18.700 ;
        RECT 12.830 14.790 13.180 18.240 ;
        RECT 13.620 15.250 13.970 18.700 ;
        RECT 14.410 14.790 14.760 18.240 ;
        RECT 15.200 15.250 15.550 18.700 ;
        RECT 15.990 14.790 16.340 18.240 ;
        RECT 6.350 13.760 16.340 14.790 ;
        RECT 8.750 11.760 9.650 13.760 ;
        RECT 16.600 11.760 17.800 12.960 ;
      LAYER via3 ;
        RECT 0.700 20.660 1.700 21.660 ;
        RECT 8.780 19.790 9.620 21.730 ;
        RECT 8.780 11.790 9.620 13.730 ;
        RECT 16.700 11.860 17.700 12.860 ;
  END
END tt_asw_1v8
END LIBRARY

