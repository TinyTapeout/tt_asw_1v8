* NGSPICE file created from tt_asw_1v8_parax.ext - technology: sky130A

.subckt tt_asw_1v8_parax VGND VPWR mod bus ctrl
X0 VPWR.t14 ctrl.t0 a_264_2813.t2 VPWR.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.5 l=0.15
**devattr s=9900,366 d=18600,724
X1 bus.t6 a_264_2813.t3 mod.t6 VPWR.t10 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=17400,658 d=17400,658
X2 a_264_2813.t0 ctrl.t1 VPWR.t12 VPWR.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.5 l=0.15
**devattr s=18600,724 d=9900,366
X3 a_680_3582# a_264_2813.t4 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.15
**devattr s=17400,716 d=17400,716
X4 bus.t10 a_680_3582# mod.t9 VGND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=17400,658 d=17400,658
X5 mod.t5 a_264_2813.t5 bus.t5 VPWR.t9 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=17400,658 d=17400,658
X6 bus.t4 a_264_2813.t6 mod.t1 VPWR.t8 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=17400,658 d=34800,1316
X7 bus.t3 a_264_2813.t7 mod.t4 VPWR.t7 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=34800,1316 d=17400,658
X8 VPWR.t6 a_264_2813.t8 a_680_3582# VPWR.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.2475 ps=1.83 w=1.5 l=0.15
**devattr s=9900,366 d=18600,724
X9 mod.t10 a_680_3582# bus.t9 VGND.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=17400,658 d=34800,1316
X10 bus.t2 a_264_2813.t9 mod.t0 VPWR.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=17400,658 d=17400,658
X11 a_264_2813.t1 ctrl.t2 VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.5 l=0.15
**devattr s=17400,716 d=17400,716
X12 bus.t8 a_680_3582# mod.t8 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=34800,1316 d=17400,658
X13 mod.t2 a_264_2813.t10 bus.t1 VPWR.t3 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=17400,658 d=17400,658
X14 a_680_3582# a_264_2813.t11 VPWR.t2 VPWR.t1 sky130_fd_pr__pfet_01v8 ad=0.2475 pd=1.83 as=0 ps=0 w=1.5 l=0.15
**devattr s=18600,724 d=9900,366
X15 mod.t3 a_264_2813.t12 bus.t0 VPWR.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=17400,658 d=17400,658
X16 mod.t7 a_680_3582# bus.t7 VGND.t4 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=3 l=0.5
**devattr s=17400,658 d=17400,658
R0 ctrl.n1 ctrl.t0 317.212
R1 ctrl.t0 ctrl.n0 317.212
R2 ctrl.n1 ctrl.t1 317.185
R3 ctrl.t1 ctrl.n0 317.185
R4 ctrl.n3 ctrl.t2 231.677
R5 ctrl.n2 ctrl.n1 68.35
R6 ctrl.n2 ctrl.n0 66.8028
R7 ctrl ctrl.n3 9.07858
R8 ctrl.n3 ctrl.n2 0.387869
R9 a_264_2813.n2 a_264_2813.t6 337.178
R10 a_264_2813.n0 a_264_2813.t6 337.178
R11 a_264_2813.n1 a_264_2813.t7 336.748
R12 a_264_2813.t7 a_264_2813.n3 336.748
R13 a_264_2813.n1 a_264_2813.t10 336.748
R14 a_264_2813.t10 a_264_2813.n3 336.748
R15 a_264_2813.t3 a_264_2813.n1 336.748
R16 a_264_2813.n3 a_264_2813.t3 336.748
R17 a_264_2813.t5 a_264_2813.n1 336.748
R18 a_264_2813.n3 a_264_2813.t5 336.748
R19 a_264_2813.n0 a_264_2813.t9 336.748
R20 a_264_2813.t9 a_264_2813.n2 336.748
R21 a_264_2813.n0 a_264_2813.t12 336.748
R22 a_264_2813.t12 a_264_2813.n2 336.748
R23 a_264_2813.n7 a_264_2813.t8 317.212
R24 a_264_2813.t8 a_264_2813.n6 317.212
R25 a_264_2813.t11 a_264_2813.n6 317.185
R26 a_264_2813.n7 a_264_2813.t11 317.185
R27 a_264_2813.n4 a_264_2813.t4 231.684
R28 a_264_2813.n9 a_264_2813.n8 150.726
R29 a_264_2813.n4 a_264_2813.n6 68.09
R30 a_264_2813.n4 a_264_2813.n7 67.0628
R31 a_264_2813.n8 a_264_2813.t1 62.2152
R32 a_264_2813.n9 a_264_2813.t2 21.6705
R33 a_264_2813.t0 a_264_2813.n9 21.6705
R34 a_264_2813.n4 a_264_2813.n5 7.113
R35 a_264_2813.n8 a_264_2813.n4 5.22455
R36 a_264_2813.n3 a_264_2813.n2 2.14724
R37 a_264_2813.n1 a_264_2813.n0 2.14724
R38 a_264_2813.n5 a_264_2813.n1 1.41083
R39 a_264_2813.n5 a_264_2813.n3 1.39452
R40 VPWR.n9 VPWR.n5 3938.82
R41 VPWR.n9 VPWR.n6 3938.82
R42 VPWR.n10 VPWR.n6 3938.82
R43 VPWR.n10 VPWR.n5 3938.82
R44 VPWR.n30 VPWR.n15 1796.47
R45 VPWR.n23 VPWR.n22 1796.47
R46 VPWR.n22 VPWR.n19 1796.47
R47 VPWR.n32 VPWR.n15 1796.47
R48 VPWR.n26 VPWR.n17 1055.29
R49 VPWR.n26 VPWR.n16 1055.29
R50 VPWR.n30 VPWR.n17 741.178
R51 VPWR.n23 VPWR.n17 741.178
R52 VPWR.n32 VPWR.n16 741.178
R53 VPWR.n19 VPWR.n16 741.178
R54 VPWR.n8 VPWR.n7 420.142
R55 VPWR.n8 VPWR.n4 420.142
R56 VPWR.t5 VPWR.n15 234.965
R57 VPWR.n22 VPWR.t11 234.965
R58 VPWR.n25 VPWR.t1 208.537
R59 VPWR.n25 VPWR.t13 208.537
R60 VPWR.t8 VPWR.n5 193.457
R61 VPWR.t7 VPWR.n6 193.457
R62 VPWR.n21 VPWR.n18 191.625
R63 VPWR.n29 VPWR.n13 191.625
R64 VPWR.n1 VPWR.t12 174.149
R65 VPWR.n1 VPWR.t14 174.053
R66 VPWR.n2 VPWR.t2 174.053
R67 VPWR.n3 VPWR.t6 174.053
R68 VPWR.n7 VPWR.n0 169.036
R69 VPWR.n12 VPWR.n4 169.036
R70 VPWR.t0 VPWR.t8 144.606
R71 VPWR.t4 VPWR.t0 144.606
R72 VPWR.t9 VPWR.t4 144.606
R73 VPWR.t9 VPWR.t10 144.606
R74 VPWR.t10 VPWR.t3 144.606
R75 VPWR.t3 VPWR.t7 144.606
R76 VPWR.n21 VPWR.n20 132.25
R77 VPWR.n34 VPWR.n13 112.566
R78 VPWR.n28 VPWR.n27 112.566
R79 VPWR.n27 VPWR.n14 112.566
R80 VPWR.n29 VPWR.n28 79.0593
R81 VPWR.n28 VPWR.n18 79.0593
R82 VPWR.n31 VPWR.t5 61.7891
R83 VPWR.n31 VPWR.t1 61.7891
R84 VPWR.t13 VPWR.n24 61.7891
R85 VPWR.n24 VPWR.t11 61.7891
R86 VPWR.n30 VPWR.n29 46.2505
R87 VPWR.n31 VPWR.n30 46.2505
R88 VPWR.n23 VPWR.n18 46.2505
R89 VPWR.n24 VPWR.n23 46.2505
R90 VPWR.n20 VPWR.n19 46.2505
R91 VPWR.n24 VPWR.n19 46.2505
R92 VPWR.n33 VPWR.n32 46.2505
R93 VPWR.n32 VPWR.n31 46.2505
R94 VPWR.n35 VPWR.n34 32.1236
R95 VPWR.n22 VPWR.n21 26.4291
R96 VPWR.n15 VPWR.n13 26.4291
R97 VPWR.n27 VPWR.n26 26.4291
R98 VPWR.n26 VPWR.n25 26.4291
R99 VPWR.n7 VPWR.n5 16.8187
R100 VPWR.n6 VPWR.n4 16.8187
R101 VPWR.n11 VPWR.n0 15.5801
R102 VPWR.n12 VPWR.n11 15.5801
R103 VPWR.n35 VPWR.n12 12.1309
R104 VPWR.n9 VPWR.n8 10.8829
R105 VPWR.t9 VPWR.n9 10.8829
R106 VPWR.n11 VPWR.n10 10.8829
R107 VPWR.n10 VPWR.t9 10.8829
R108 VPWR.n34 VPWR.n33 8.61589
R109 VPWR.n33 VPWR.n14 8.61589
R110 VPWR.n20 VPWR.n14 8.61589
R111 VPWR.n37 VPWR.n0 4.54886
R112 VPWR.n38 VPWR.n37 2.2055
R113 VPWR.n37 VPWR.n36 0.901542
R114 VPWR.n38 VPWR 0.4846
R115 VPWR.n36 VPWR.n3 0.46925
R116 VPWR VPWR.n38 0.368667
R117 VPWR.n36 VPWR.n35 0.211864
R118 VPWR.n2 VPWR.n1 0.122375
R119 VPWR.n3 VPWR.n2 0.097375
R120 mod.n5 mod.t4 85.0593
R121 mod.n3 mod.n2 75.6077
R122 mod.n4 mod.n0 75.5377
R123 mod.n3 mod.n1 75.5377
R124 mod.n7 mod.t8 31.41
R125 mod.n8 mod.t10 31.34
R126 mod.n7 mod.n6 25.54
R127 mod.n0 mod.t6 9.52217
R128 mod.n0 mod.t2 9.52217
R129 mod.n1 mod.t0 9.52217
R130 mod.n1 mod.t5 9.52217
R131 mod.n2 mod.t1 9.52217
R132 mod.n2 mod.t3 9.52217
R133 mod.n6 mod.t9 5.8005
R134 mod.n6 mod.t7 5.8005
R135 mod.n10 mod.n9 0.393722
R136 mod.n4 mod.n3 0.0705566
R137 mod.n5 mod.n4 0.0705566
R138 mod.n8 mod.n7 0.0705566
R139 mod.n9 mod.n5 0.0641274
R140 mod mod.n10 0.0527222
R141 mod.n10 mod 0.0527222
R142 mod.n9 mod.n8 0.0140236
R143 bus.n3 bus.t4 85.1314
R144 bus.n3 bus.n2 75.5377
R145 bus.n4 bus.n1 75.5377
R146 bus.n5 bus.n0 75.5377
R147 bus.n8 bus.n7 25.6121
R148 bus.n8 bus.n6 25.54
R149 bus.n2 bus.t0 9.52217
R150 bus.n2 bus.t2 9.52217
R151 bus.n1 bus.t5 9.52217
R152 bus.n1 bus.t6 9.52217
R153 bus.n0 bus.t1 9.52217
R154 bus.n0 bus.t3 9.52217
R155 bus.n6 bus.t9 5.8005
R156 bus.n6 bus.t10 5.8005
R157 bus.n7 bus.t7 5.8005
R158 bus.n7 bus.t8 5.8005
R159 bus.n10 bus.n9 0.393722
R160 bus.n9 bus.n5 0.102029
R161 bus.n4 bus.n3 0.0725971
R162 bus.n5 bus.n4 0.0725971
R163 bus bus.n10 0.0527222
R164 bus.n10 bus 0.0527222
R165 bus.n9 bus.n8 0.050466
R166 VGND.n20 VGND.n19 80126.8
R167 VGND.n18 VGND.n13 5040.88
R168 VGND.n18 VGND.n14 5040.88
R169 VGND.n23 VGND.n13 5040.88
R170 VGND.n23 VGND.n14 5040.88
R171 VGND.n31 VGND.n5 2595.76
R172 VGND.n32 VGND.n5 2595.76
R173 VGND.n36 VGND.n3 2595.76
R174 VGND.n9 VGND.n4 1680.29
R175 VGND.n33 VGND.n4 1680.29
R176 VGND.t5 VGND.t4 1384.86
R177 VGND.n31 VGND.n9 915.471
R178 VGND.n9 VGND.n3 915.471
R179 VGND.n33 VGND.n32 915.471
R180 VGND.n34 VGND.n33 915.471
R181 VGND.n22 VGND.n7 905.883
R182 VGND.t6 VGND.n19 832.549
R183 VGND.n22 VGND.t5 832.549
R184 VGND.t4 VGND.n15 692.431
R185 VGND.t5 VGND.t4 681.569
R186 VGND.t0 VGND.n7 681.569
R187 VGND.t0 VGND.n8 681.569
R188 VGND.n8 VGND.t2 681.569
R189 VGND.n36 VGND.n35 543.638
R190 VGND.t7 VGND.t6 456.767
R191 VGND.t4 VGND.n21 340.784
R192 VGND.n17 VGND.n12 327.529
R193 VGND.n24 VGND.n12 327.529
R194 VGND.n34 VGND.n2 292.5
R195 VGND.n32 VGND.n6 292.5
R196 VGND.n32 VGND.t0 292.5
R197 VGND.n31 VGND.n30 292.5
R198 VGND.t0 VGND.n31 292.5
R199 VGND.n3 VGND.n1 292.5
R200 VGND.t2 VGND.n3 292.5
R201 VGND.n20 VGND.t7 208.148
R202 VGND.n35 VGND.n34 207.823
R203 VGND.n37 VGND.n2 168.66
R204 VGND.n10 VGND.n6 168.66
R205 VGND.n17 VGND.n16 165.648
R206 VGND.n25 VGND.n24 165.648
R207 VGND.n38 VGND.n37 110.314
R208 VGND.n28 VGND.n27 109.177
R209 VGND.n29 VGND.n28 108.424
R210 VGND.n26 VGND.n10 108.424
R211 VGND.n28 VGND.n4 83.5719
R212 VGND.n8 VGND.n4 83.5719
R213 VGND.n37 VGND.n36 83.5719
R214 VGND.n10 VGND.n5 83.5719
R215 VGND.n7 VGND.n5 83.5719
R216 VGND.n0 VGND.t1 64.0037
R217 VGND.n40 VGND.t3 62.2777
R218 VGND.n20 VGND.n15 61.3551
R219 VGND.n35 VGND.t2 61.2599
R220 VGND.n27 VGND.n6 59.4829
R221 VGND.n27 VGND.n2 59.4829
R222 VGND.n14 VGND.n12 58.5005
R223 VGND.n15 VGND.n14 58.5005
R224 VGND.n13 VGND.n11 58.5005
R225 VGND.n21 VGND.n13 58.5005
R226 VGND.n24 VGND.n23 53.1823
R227 VGND.n23 VGND.n22 53.1823
R228 VGND.n18 VGND.n17 53.1823
R229 VGND.n19 VGND.n18 53.1823
R230 VGND.n21 VGND.n20 30.1966
R231 VGND.n16 VGND.n11 9.79409
R232 VGND.n25 VGND.n11 9.79409
R233 VGND.n26 VGND.n25 7.82865
R234 VGND.n30 VGND.n26 6.09207
R235 VGND.n30 VGND.n29 6.09207
R236 VGND.n29 VGND.n1 6.09207
R237 VGND.n38 VGND.n1 4.20291
R238 VGND.n16 VGND.n0 3.61335
R239 VGND.n41 VGND.n40 1.7055
R240 VGND.n39 VGND.n38 1.03383
R241 VGND.n41 VGND 0.829267
R242 VGND.n40 VGND.n39 0.5005
R243 VGND.n39 VGND.n0 0.2005
R244 VGND VGND.n41 0.024
C0 a_680_3582# bus 0.373525f
C1 ctrl bus 0.002912f
C2 a_680_3582# mod 0.821024f
C3 bus VPWR 1.31714f
C4 ctrl mod 0.23001f
C5 mod VPWR 0.471489f
C6 ctrl a_680_3582# 0.130281f
C7 a_680_3582# VPWR 0.863753f
C8 ctrl VPWR 1.06756f
C9 bus mod 8.507401f
.ends

