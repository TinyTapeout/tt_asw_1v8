magic
tech sky130A
magscale 1 2
timestamp 1711041971
<< pwell >>
rect 970 3450 1060 3510
rect 2380 2690 2810 2750
<< psubdiff >>
rect 462 1416 614 1440
rect 462 1222 614 1246
<< psubdiffcont >>
rect 462 1246 614 1416
<< locali >>
rect 462 1416 614 1432
rect 462 1230 614 1246
<< viali >>
rect 1546 3356 1594 3404
rect 2836 3126 2884 3174
rect 1546 2156 1594 2204
<< metal1 >>
rect 2254 4130 2260 4210
rect 2340 4130 3290 4210
rect 684 3970 690 4030
rect 750 3970 756 4030
rect 690 3915 1440 3970
rect 1668 3915 1674 3916
rect 690 3910 1674 3915
rect 690 3740 750 3910
rect 1375 3865 1674 3910
rect 1380 3750 1440 3865
rect 1668 3864 1674 3865
rect 1726 3864 1732 3916
rect 1880 3860 3040 3920
rect 415 3451 421 3510
rect 480 3451 689 3510
rect 730 3450 1290 3510
rect 1430 3450 1780 3510
rect 1840 3450 1846 3510
rect 680 2970 740 3180
rect 674 2910 680 2970
rect 740 2910 746 2970
rect 970 2940 1030 3450
rect 1710 3410 1770 3450
rect 1534 3404 1770 3410
rect 1534 3356 1546 3404
rect 1594 3356 1770 3404
rect 1534 3350 1770 3356
rect 1674 3181 1726 3187
rect 1280 3130 1674 3180
rect 1674 3123 1726 3129
rect 1880 2940 1940 3860
rect 2226 3690 2236 3746
rect 2296 3690 2306 3746
rect 2418 3692 2428 3748
rect 2488 3692 2498 3748
rect 2610 3692 2620 3748
rect 2680 3692 2690 3748
rect 2806 3688 2816 3744
rect 2876 3688 2886 3744
rect 2996 3692 3006 3748
rect 3066 3692 3076 3748
rect 3210 3560 3290 4130
rect 2324 3492 2334 3548
rect 2394 3492 2404 3548
rect 2512 3494 2522 3550
rect 2582 3494 2592 3550
rect 2710 3492 2720 3548
rect 2780 3492 2790 3548
rect 2898 3488 2908 3544
rect 2968 3488 2978 3544
rect 3114 3480 3120 3560
rect 3200 3480 3290 3560
rect 2280 3220 2940 3280
rect 2380 2940 2440 3220
rect 2830 3174 2890 3186
rect 2830 3126 2836 3174
rect 2884 3126 2890 3174
rect 2830 3040 2890 3126
rect 2970 3040 3030 3046
rect 2830 2980 2970 3040
rect 2970 2974 3030 2980
rect 970 2880 2440 2940
rect 538 2644 544 2696
rect 596 2695 602 2696
rect 596 2690 795 2695
rect 970 2690 1030 2880
rect 1650 2690 1710 2696
rect 2380 2690 2880 2750
rect 596 2645 1650 2690
rect 596 2644 602 2645
rect 690 2630 1650 2645
rect 380 2560 440 2566
rect 380 2090 440 2500
rect 690 2340 740 2630
rect 1390 2360 1440 2630
rect 1650 2624 1710 2630
rect 2326 2398 2336 2452
rect 2388 2398 2398 2452
rect 2520 2398 2530 2452
rect 2582 2398 2592 2452
rect 2232 2244 2242 2298
rect 2294 2244 2304 2298
rect 2422 2244 2432 2298
rect 2484 2244 2494 2298
rect 2618 2242 2628 2296
rect 2680 2242 2690 2296
rect 1534 2204 1800 2210
rect 1534 2156 1546 2204
rect 1594 2156 1800 2204
rect 1534 2150 1800 2156
rect 1740 2090 1800 2150
rect 380 2030 690 2090
rect 730 2030 1290 2090
rect 1440 2030 1800 2090
rect 2280 2060 2540 2120
rect 970 1900 1030 2030
rect 964 1840 970 1900
rect 1030 1840 1036 1900
rect 1740 1790 1800 2030
rect 2380 1920 2440 2060
rect 2380 1854 2440 1860
rect 2600 1920 2660 1926
rect 2820 1920 2880 2690
rect 3210 2310 3290 3480
rect 3064 2230 3070 2310
rect 3150 2230 3290 2310
rect 2660 1860 2880 1920
rect 2600 1854 2660 1860
rect 538 1524 544 1576
rect 596 1575 602 1576
rect 690 1575 740 1780
rect 596 1525 740 1575
rect 596 1524 602 1525
rect 690 1520 740 1525
rect 463 1359 622 1439
rect 1280 1420 1340 1780
rect 1740 1730 3070 1790
rect 3130 1730 3136 1790
rect 1650 1670 1710 1676
rect 1650 1420 1710 1610
rect 1280 1360 1710 1420
rect 457 1200 463 1359
rect 622 1200 628 1359
<< via1 >>
rect 2260 4130 2340 4210
rect 690 3970 750 4030
rect 1674 3864 1726 3916
rect 421 3451 480 3510
rect 1780 3450 1840 3510
rect 680 2910 740 2970
rect 1674 3129 1726 3181
rect 2236 3690 2296 3746
rect 2428 3692 2488 3748
rect 2620 3692 2680 3748
rect 2816 3688 2876 3744
rect 3006 3692 3066 3748
rect 2334 3492 2394 3548
rect 2522 3494 2582 3550
rect 2720 3492 2780 3548
rect 2908 3488 2968 3544
rect 3120 3480 3200 3560
rect 2970 2980 3030 3040
rect 544 2644 596 2696
rect 1650 2630 1710 2690
rect 380 2500 440 2560
rect 2336 2398 2388 2452
rect 2530 2398 2582 2452
rect 2242 2244 2294 2298
rect 2432 2244 2484 2298
rect 2628 2242 2680 2296
rect 970 1840 1030 1900
rect 2380 1860 2440 1920
rect 3070 2230 3150 2310
rect 2600 1860 2660 1920
rect 544 1524 596 1576
rect 3070 1730 3130 1790
rect 1650 1610 1710 1670
rect 463 1200 622 1359
<< metal2 >>
rect 2260 4210 2340 4216
rect 690 4140 750 4149
rect 2011 4130 2020 4210
rect 2100 4130 2260 4210
rect 2260 4124 2340 4130
rect 690 4030 750 4080
rect 750 3970 930 4030
rect 690 3964 750 3970
rect 272 3451 281 3511
rect 341 3510 350 3511
rect 421 3510 480 3516
rect 341 3451 421 3510
rect 421 3445 480 3451
rect 680 2970 740 2976
rect 870 2970 930 3970
rect 1674 3916 1726 3922
rect 1674 3858 1726 3864
rect 1675 3181 1725 3858
rect 2236 3755 2296 3756
rect 2428 3755 2488 3758
rect 2620 3755 2680 3758
rect 3006 3755 3066 3758
rect 2015 3748 3085 3755
rect 2015 3746 2428 3748
rect 2015 3690 2236 3746
rect 2296 3692 2428 3746
rect 2488 3692 2620 3748
rect 2680 3744 3006 3748
rect 2680 3692 2816 3744
rect 2296 3690 2816 3692
rect 2015 3688 2816 3690
rect 2876 3692 3006 3744
rect 3066 3692 3085 3748
rect 2876 3688 3085 3692
rect 2015 3685 3085 3688
rect 1780 3510 1840 3516
rect 1840 3450 1880 3510
rect 1940 3450 1949 3510
rect 1780 3444 1840 3450
rect 1668 3129 1674 3181
rect 1726 3129 1732 3181
rect 740 2910 930 2970
rect 680 2904 740 2910
rect 544 2696 596 2702
rect 544 2638 596 2644
rect 211 2500 220 2560
rect 280 2500 380 2560
rect 440 2500 446 2560
rect 545 1582 595 2638
rect 1644 2630 1650 2690
rect 1710 2630 1716 2690
rect 970 1900 1030 1906
rect 544 1576 596 1582
rect 544 1518 596 1524
rect 970 1560 1030 1840
rect 1650 1670 1710 2630
rect 2015 2615 2085 3685
rect 2236 3680 2296 3685
rect 2428 3682 2488 3685
rect 2620 3682 2680 3685
rect 2816 3678 2876 3685
rect 3006 3682 3066 3685
rect 3120 3560 3200 3566
rect 2220 3550 3120 3560
rect 2220 3548 2522 3550
rect 2220 3492 2334 3548
rect 2394 3494 2522 3548
rect 2582 3548 3120 3550
rect 2582 3494 2720 3548
rect 2394 3492 2720 3494
rect 2780 3544 3120 3548
rect 2780 3492 2908 3544
rect 2220 3488 2908 3492
rect 2968 3488 3120 3544
rect 2220 3480 3120 3488
rect 2908 3478 2968 3480
rect 3120 3474 3200 3480
rect 3122 3040 3178 3047
rect 2964 2980 2970 3040
rect 3030 3038 3180 3040
rect 3030 2982 3122 3038
rect 3178 2982 3180 3038
rect 3030 2980 3180 2982
rect 3122 2973 3178 2980
rect 2006 2545 2015 2615
rect 2085 2545 2094 2615
rect 2015 2460 2085 2545
rect 2336 2460 2388 2462
rect 2530 2460 2582 2462
rect 2009 2452 2675 2460
rect 2009 2398 2336 2452
rect 2388 2398 2530 2452
rect 2582 2398 2675 2452
rect 2009 2390 2675 2398
rect 2336 2388 2388 2390
rect 2530 2388 2582 2390
rect 3070 2310 3150 2316
rect 2140 2298 3070 2310
rect 2140 2244 2242 2298
rect 2294 2244 2432 2298
rect 2484 2296 3070 2298
rect 2484 2244 2628 2296
rect 2140 2242 2628 2244
rect 2680 2242 3070 2296
rect 2140 2230 3070 2242
rect 3070 2224 3150 2230
rect 2374 1860 2380 1920
rect 2440 1860 2600 1920
rect 2660 1860 2666 1920
rect 1644 1610 1650 1670
rect 1710 1610 1716 1670
rect 2380 1560 2440 1860
rect 3070 1790 3130 1796
rect 3130 1730 3200 1790
rect 3260 1730 3269 1790
rect 3070 1724 3130 1730
rect 970 1500 2440 1560
rect 463 1359 622 1365
rect 463 1147 622 1200
rect 458 998 467 1147
rect 617 998 626 1147
rect 463 993 622 998
<< via2 >>
rect 690 4080 750 4140
rect 2020 4130 2100 4210
rect 281 3451 341 3511
rect 1880 3450 1940 3510
rect 220 2500 280 2560
rect 3122 2982 3178 3038
rect 2015 2545 2085 2615
rect 3200 1730 3260 1790
rect 467 998 617 1147
<< metal3 >>
rect 120 4346 360 4352
rect 120 2358 126 4346
rect 354 2358 360 4346
rect 890 4300 950 4352
rect 690 4240 950 4300
rect 690 4145 750 4240
rect 685 4140 755 4145
rect 685 4080 690 4140
rect 750 4080 755 4140
rect 890 4130 950 4240
rect 1750 4346 1930 4352
rect 685 4075 755 4080
rect 1750 3958 1756 4346
rect 1924 4210 1930 4346
rect 3320 4346 3560 4352
rect 2015 4210 2105 4215
rect 1924 4130 2020 4210
rect 2100 4130 2105 4210
rect 1924 3958 1930 4130
rect 2015 4125 2105 4130
rect 1750 3952 1930 3958
rect 1875 3510 1945 3515
rect 3320 3510 3326 4346
rect 1875 3450 1880 3510
rect 1940 3450 3326 3510
rect 1875 3445 1945 3450
rect 3117 3040 3183 3043
rect 3320 3040 3326 3450
rect 3117 3038 3326 3040
rect 3117 2982 3122 3038
rect 3178 2982 3326 3038
rect 3117 2980 3326 2982
rect 3117 2977 3183 2980
rect 120 2352 360 2358
rect 1750 2746 1930 2752
rect 1750 2358 1756 2746
rect 1924 2615 1930 2746
rect 2010 2615 2090 2620
rect 1924 2545 2015 2615
rect 2085 2545 2090 2615
rect 1924 2358 1930 2545
rect 2010 2540 2090 2545
rect 1750 2352 1930 2358
rect 3320 2358 3326 2980
rect 3554 2358 3560 4346
rect 3320 2352 3560 2358
rect 3195 1790 3265 1795
rect 3372 1790 3378 1792
rect 3195 1730 3200 1790
rect 3260 1730 3378 1790
rect 3195 1725 3265 1730
rect 3372 1728 3378 1730
rect 3442 1728 3448 1792
rect 462 1147 622 1152
rect 462 1027 467 1147
rect 423 1021 467 1027
rect 617 1027 622 1147
rect 617 1021 661 1027
rect 423 777 661 783
<< via3 >>
rect 126 3511 354 4346
rect 126 3451 281 3511
rect 281 3451 341 3511
rect 341 3451 354 3511
rect 126 2560 354 3451
rect 126 2500 220 2560
rect 220 2500 280 2560
rect 280 2500 354 2560
rect 126 2358 354 2500
rect 1756 3958 1924 4346
rect 1756 2358 1924 2746
rect 3326 2358 3554 4346
rect 3378 1728 3442 1792
rect 423 998 467 1021
rect 467 998 617 1021
rect 617 998 661 1021
rect 423 783 661 998
<< metal4 >>
rect 120 4346 360 4352
rect 120 2358 126 4346
rect 354 2358 360 4346
rect 1750 4346 1930 4352
rect 1750 3958 1756 4346
rect 1924 3958 1930 4346
rect 1750 3952 1930 3958
rect 3320 4346 3560 4352
rect 120 1022 360 2358
rect 1750 2746 1930 2752
rect 1750 2358 1756 2746
rect 1924 2358 1930 2746
rect 1750 2352 1930 2358
rect 3320 2358 3326 4346
rect 3554 2358 3560 4346
rect 3320 1792 3560 2358
rect 3320 1728 3378 1792
rect 3442 1728 3560 1792
rect 120 1021 662 1022
rect 120 783 423 1021
rect 661 783 662 1021
rect 120 782 662 783
rect 120 0 360 782
rect 3320 0 3560 1728
use sky130_fd_pr__nfet_01v8_H7HSAV  XM1
timestamp 1711022820
transform 1 0 711 0 1 3460
box -211 -460 211 460
use sky130_fd_pr__pfet_01v8_XJT9DL  XM2
timestamp 1711022820
transform 1 0 1363 0 1 3469
box -263 -469 263 469
use sky130_fd_pr__nfet_01v8_5ZNSAF  XM3
timestamp 1711022820
transform 1 0 2459 0 1 2400
box -359 -460 359 460
use sky130_fd_pr__pfet_01v8_XJT9DL  XM4
timestamp 1711022820
transform 1 0 1363 0 1 2069
box -263 -469 263 469
use sky130_fd_pr__pfet_01v8_XJKGNP  XM4A
timestamp 1711022820
transform 1 0 2651 0 1 3569
box -551 -469 551 469
use sky130_fd_pr__nfet_01v8_H7HSAV  XM5
timestamp 1711022820
transform 1 0 711 0 1 2060
box -211 -460 211 460
<< labels >>
rlabel metal4 3320 0 3560 4352 1 VPWR
port 2 n power input
rlabel metal4 1750 3952 1930 4352 1 mod
port 3 n analog bidirectional
rlabel metal4 1750 2352 1930 2752 1 bus
port 4 n analog bidirectional
rlabel metal3 890 4172 950 4352 1 ctrl
port 5 n signal input
rlabel metal4 120 0 360 4352 1 VGND
port 1 n ground input
flabel metal1 970 2640 1030 3500 0 FreeSans 160 0 0 0 tgon_n
flabel metal1 730 2030 1290 2090 0 FreeSans 160 0 0 0 tgon
<< properties >>
string FIXED_BBOX 0 0 3680 4352
<< end >>
