magic
tech sky130A
magscale 1 2
timestamp 1711022820
<< error_p >>
rect 19 331 77 337
rect 19 297 31 331
rect 19 291 77 297
rect -77 -297 -19 -291
rect -77 -331 -65 -297
rect -77 -337 -19 -331
<< nwell >>
rect -263 -469 263 469
<< pmos >>
rect -63 -250 -33 250
rect 33 -250 63 250
<< pdiff >>
rect -125 238 -63 250
rect -125 -238 -113 238
rect -79 -238 -63 238
rect -125 -250 -63 -238
rect -33 238 33 250
rect -33 -238 -17 238
rect 17 -238 33 238
rect -33 -250 33 -238
rect 63 238 125 250
rect 63 -238 79 238
rect 113 -238 125 238
rect 63 -250 125 -238
<< pdiffc >>
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
<< nsubdiff >>
rect -227 399 -131 433
rect 131 399 227 433
rect -227 337 -193 399
rect 193 337 227 399
rect -227 -399 -193 -337
rect 193 -399 227 -337
rect -227 -433 -131 -399
rect 131 -433 227 -399
<< nsubdiffcont >>
rect -131 399 131 433
rect -227 -337 -193 337
rect 193 -337 227 337
rect -131 -433 131 -399
<< poly >>
rect 15 331 81 347
rect 15 297 31 331
rect 65 297 81 331
rect 15 281 81 297
rect -63 250 -33 276
rect 33 250 63 281
rect -63 -281 -33 -250
rect 33 -276 63 -250
rect -81 -297 -15 -281
rect -81 -331 -65 -297
rect -31 -331 -15 -297
rect -81 -347 -15 -331
<< polycont >>
rect 31 297 65 331
rect -65 -331 -31 -297
<< locali >>
rect -227 399 -131 433
rect 131 399 227 433
rect -227 337 -193 399
rect 193 337 227 399
rect 15 297 31 331
rect 65 297 81 331
rect -113 238 -79 254
rect -113 -254 -79 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 79 238 113 254
rect 79 -254 113 -238
rect -81 -331 -65 -297
rect -31 -331 -15 -297
rect -227 -399 -193 -337
rect 193 -399 227 -337
rect -227 -433 -131 -399
rect 131 -433 227 -399
<< viali >>
rect 31 297 65 331
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
rect -65 -331 -31 -297
<< metal1 >>
rect 19 331 77 337
rect 19 297 31 331
rect 65 297 77 331
rect 19 291 77 297
rect -119 238 -73 250
rect -119 -238 -113 238
rect -79 -238 -73 238
rect -119 -250 -73 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 73 238 119 250
rect 73 -238 79 238
rect 113 -238 119 238
rect 73 -250 119 -238
rect -77 -297 -19 -291
rect -77 -331 -65 -297
rect -31 -331 -19 -297
rect -77 -337 -19 -331
<< properties >>
string FIXED_BBOX -210 -416 210 416
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
