* NGSPICE file created from tt_asw_1v8_parax.ext - technology: sky130A

.subckt tt_asw_1v8_parax VGND VPWR mod bus ctrl
X0 bus.t10 a_726_1810# mod.t10 VGND.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=16500,566
X1 mod.t0 tgon_n.t3 bus.t0 VPWR.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=16500,566
X2 tgon_n.t1 ctrl.t0 VPWR.t13 VPWR.t12 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=31000,1124
X3 a_726_1810# tgon_n.t4 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0 ps=0 w=2.5 l=0.15
**devattr s=29000,1116 d=29000,1116
X4 mod.t7 a_726_1810# bus.t9 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=16500,566
X5 VPWR.t15 ctrl.t1 tgon_n.t2 VPWR.t14 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=31000,1124 d=16500,566
X6 a_726_1810# tgon_n.t5 VPWR.t10 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.775 pd=5.62 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=31000,1124
X7 mod.t11 tgon_n.t6 bus.t11 VPWR.t8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=16500,566
X8 bus.t8 a_726_1810# mod.t8 VGND.t3 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=31000,1124 d=16500,566
X9 bus.t4 tgon_n.t7 mod.t4 VPWR.t7 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=16500,566
X10 VPWR.t6 tgon_n.t8 a_726_1810# VPWR.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.775 ps=5.62 w=2.5 l=0.15
**devattr s=31000,1124 d=16500,566
X11 mod.t9 a_726_1810# bus.t7 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=31000,1124
X12 bus.t6 tgon_n.t9 mod.t6 VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=16500,566
X13 mod.t1 tgon_n.t10 bus.t1 VPWR.t3 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=16500,566
X14 bus.t3 tgon_n.t11 mod.t3 VPWR.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=31000,1124
X15 mod.t2 tgon_n.t12 bus.t2 VPWR.t1 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=31000,1124 d=16500,566
X16 tgon_n.t0 ctrl.t2 VGND.t6 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=29000,1116 d=29000,1116
X17 bus.t5 tgon_n.t13 mod.t5 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.5 l=0.15
**devattr s=16500,566 d=16500,566
R0 mod.n5 mod.n3 89.7951
R1 mod.n9 mod.n8 89.5122
R2 mod.n7 mod.n6 89.5013
R3 mod.n5 mod.n4 89.4959
R4 mod.n1 mod.t8 40.7986
R5 mod.n2 mod.t9 40.5071
R6 mod.n1 mod.n0 32.5817
R7 mod.n3 mod.t6 13.0025
R8 mod.n3 mod.t2 13.0025
R9 mod.n4 mod.t5 13.0025
R10 mod.n4 mod.t11 13.0025
R11 mod.n6 mod.t4 13.0025
R12 mod.n6 mod.t1 13.0025
R13 mod.n8 mod.t3 13.0025
R14 mod.n8 mod.t0 13.0025
R15 mod.n11 mod.n10 11.0855
R16 mod.n0 mod.t10 7.9205
R17 mod.n0 mod.t7 7.9205
R18 mod.n10 mod.n2 7.25988
R19 mod.n10 mod.n9 4.988
R20 mod.n7 mod.n5 0.309875
R21 mod.n2 mod.n1 0.30675
R22 mod.n9 mod.n7 0.29425
R23 mod mod.n11 0.0527222
R24 mod.n11 mod 0.0527222
R25 bus.n1 bus.t3 103.12
R26 bus.n6 bus.t2 102.775
R27 bus.n5 bus.n4 89.7785
R28 bus.n3 bus.n2 89.7785
R29 bus.n1 bus.n0 89.7676
R30 bus.n9 bus.n7 32.6475
R31 bus.n9 bus.n8 32.301
R32 bus.n4 bus.t11 13.0025
R33 bus.n4 bus.t6 13.0025
R34 bus.n2 bus.t1 13.0025
R35 bus.n2 bus.t5 13.0025
R36 bus.n0 bus.t0 13.0025
R37 bus.n0 bus.t4 13.0025
R38 bus.n8 bus.t9 7.9205
R39 bus.n8 bus.t8 7.9205
R40 bus.n7 bus.t7 7.9205
R41 bus.n7 bus.t10 7.9205
R42 bus.n11 bus.n10 3.83929
R43 bus.n10 bus.n6 2.34664
R44 bus.n10 bus.n9 0.759145
R45 bus.n3 bus.n1 0.3505
R46 bus.n5 bus.n3 0.343357
R47 bus.n6 bus.n5 0.343357
R48 bus bus.n11 0.0527222
R49 bus.n11 bus 0.0527222
R50 VGND.n18 VGND.n7 33476.2
R51 VGND.n12 VGND.n8 4032.71
R52 VGND.n16 VGND.n8 4032.71
R53 VGND.n12 VGND.n10 4032.71
R54 VGND.n16 VGND.n10 4032.71
R55 VGND.n27 VGND.n4 3175.18
R56 VGND.n31 VGND.n4 3175.18
R57 VGND.n27 VGND.n5 3175.18
R58 VGND.n31 VGND.n5 3175.18
R59 VGND.n25 VGND.n19 3175.18
R60 VGND.n19 VGND.n3 3175.18
R61 VGND.n25 VGND.n20 3175.18
R62 VGND.n20 VGND.n3 3175.18
R63 VGND.n18 VGND.n17 1256.47
R64 VGND.n26 VGND.n18 720.436
R65 VGND.n23 VGND.n20 292.5
R66 VGND.n20 VGND.t0 292.5
R67 VGND.n21 VGND.n19 292.5
R68 VGND.n19 VGND.t0 292.5
R69 VGND.n29 VGND.n5 292.5
R70 VGND.n5 VGND.t0 292.5
R71 VGND.n6 VGND.n4 292.5
R72 VGND.n4 VGND.t0 292.5
R73 VGND.n13 VGND.n11 262.024
R74 VGND.n15 VGND.n11 262.024
R75 VGND.n14 VGND.n13 262.024
R76 VGND.n15 VGND.n14 262.024
R77 VGND.t2 VGND.n7 229.935
R78 VGND.n17 VGND.t3 229.935
R79 VGND.n33 VGND.n32 215.766
R80 VGND.n28 VGND.n6 206.306
R81 VGND.n30 VGND.n6 206.306
R82 VGND.n29 VGND.n28 206.306
R83 VGND.n30 VGND.n29 206.306
R84 VGND.n24 VGND.n21 206.306
R85 VGND.n22 VGND.n21 206.306
R86 VGND.n24 VGND.n23 206.306
R87 VGND.n23 VGND.n22 206.306
R88 VGND.n26 VGND.t0 159.744
R89 VGND.n32 VGND.t0 159.744
R90 VGND.t5 VGND.t2 136.258
R91 VGND.t4 VGND.t3 136.258
R92 VGND.n14 VGND.n10 83.5719
R93 VGND.n10 VGND.n9 83.5719
R94 VGND.n11 VGND.n8 83.5719
R95 VGND.n9 VGND.n8 83.5719
R96 VGND.n9 VGND.t5 68.1295
R97 VGND.n9 VGND.t4 68.1295
R98 VGND.n16 VGND.n15 58.5005
R99 VGND.n17 VGND.n16 58.5005
R100 VGND.n13 VGND.n12 58.5005
R101 VGND.n12 VGND.n7 58.5005
R102 VGND.n22 VGND.n3 58.5005
R103 VGND.n32 VGND.n3 58.5005
R104 VGND.n25 VGND.n24 58.5005
R105 VGND.n26 VGND.n25 58.5005
R106 VGND.n31 VGND.n30 58.5005
R107 VGND.n32 VGND.n31 58.5005
R108 VGND.n28 VGND.n27 58.5005
R109 VGND.n27 VGND.n26 58.5005
R110 VGND.n0 VGND.t1 44.574
R111 VGND.n0 VGND.t6 43.4058
R112 VGND VGND.n34 0.699625
R113 VGND.n2 VGND.n1 0.456792
R114 VGND.n2 VGND 0.289264
R115 VGND.n2 VGND 0.200642
R116 VGND.n1 VGND 0.196333
R117 VGND.n34 VGND 0.153642
R118 VGND.n34 VGND 0.0683118
R119 VGND.n1 VGND.n0 0.0459667
R120 VGND.n33 VGND.n2 0.0109059
R121 VGND.n34 VGND.n33 0.0109059
R122 tgon_n.n4 tgon_n.t8 650.457
R123 tgon_n.n4 tgon_n.t5 637.491
R124 tgon_n.n2 tgon_n.t3 637.274
R125 tgon_n.n0 tgon_n.t11 637.274
R126 tgon_n.n3 tgon_n.t12 637.072
R127 tgon_n.n3 tgon_n.t6 636.874
R128 tgon_n.n2 tgon_n.t10 636.874
R129 tgon_n.n1 tgon_n.t9 636.874
R130 tgon_n.n1 tgon_n.t13 636.874
R131 tgon_n.n0 tgon_n.t7 636.874
R132 tgon_n tgon_n.t4 315.099
R133 tgon_n.n6 tgon_n.t1 103.031
R134 tgon_n.n6 tgon_n.t2 102.632
R135 tgon_n tgon_n.t0 34.7176
R136 tgon_n tgon_n.n6 5.08274
R137 tgon_n.n5 tgon_n.n1 2.96092
R138 tgon_n tgon_n.n5 1.89633
R139 tgon_n.n5 tgon_n.n3 1.6255
R140 tgon_n tgon_n.n4 0.865083
R141 tgon_n.n1 tgon_n.n0 0.8005
R142 tgon_n.n3 tgon_n.n2 0.602583
R143 VPWR.n30 VPWR.n27 3165.88
R144 VPWR.n32 VPWR.n27 3165.88
R145 VPWR.n30 VPWR.n28 3165.88
R146 VPWR.n32 VPWR.n28 3165.88
R147 VPWR.n18 VPWR.n15 2149.41
R148 VPWR.n18 VPWR.n16 2149.41
R149 VPWR.n20 VPWR.n16 2149.41
R150 VPWR.n20 VPWR.n15 2149.41
R151 VPWR.n5 VPWR.n2 2149.41
R152 VPWR.n5 VPWR.n3 2149.41
R153 VPWR.n7 VPWR.n3 2149.41
R154 VPWR.n7 VPWR.n2 2149.41
R155 VPWR.n33 VPWR.n26 337.695
R156 VPWR.n29 VPWR.n26 337.695
R157 VPWR.n29 VPWR.n25 337.695
R158 VPWR.n34 VPWR.n25 256.377
R159 VPWR.n17 VPWR.n13 229.272
R160 VPWR.n17 VPWR.n14 229.272
R161 VPWR.n21 VPWR.n14 229.272
R162 VPWR.n4 VPWR.n0 229.272
R163 VPWR.n4 VPWR.n1 229.272
R164 VPWR.n8 VPWR.n1 229.272
R165 VPWR.n22 VPWR.n21 193.13
R166 VPWR.n9 VPWR.n0 184.847
R167 VPWR.t2 VPWR.n27 182.572
R168 VPWR.t1 VPWR.n28 182.572
R169 VPWR.t12 VPWR.n15 182.572
R170 VPWR.t14 VPWR.n16 182.572
R171 VPWR.n7 VPWR.t9 182.572
R172 VPWR.t5 VPWR.n5 182.572
R173 VPWR.t11 VPWR.t2 97.2286
R174 VPWR.t7 VPWR.t11 97.2286
R175 VPWR.t3 VPWR.t7 97.2286
R176 VPWR.t0 VPWR.t8 97.2286
R177 VPWR.t8 VPWR.t4 97.2286
R178 VPWR.t4 VPWR.t1 97.2286
R179 VPWR.n11 VPWR.n10 95.2965
R180 VPWR.n24 VPWR.n23 94.7212
R181 VPWR.n34 VPWR.n33 76.0476
R182 VPWR.n31 VPWR.t3 48.6146
R183 VPWR.n31 VPWR.t0 48.6146
R184 VPWR.n19 VPWR.t12 48.6146
R185 VPWR.n19 VPWR.t14 48.6146
R186 VPWR.t9 VPWR.n6 48.6146
R187 VPWR.n6 VPWR.t5 48.6146
R188 VPWR.n18 VPWR.n17 46.2505
R189 VPWR.n19 VPWR.n18 46.2505
R190 VPWR.n21 VPWR.n20 46.2505
R191 VPWR.n20 VPWR.n19 46.2505
R192 VPWR.n2 VPWR.n0 46.2505
R193 VPWR.n6 VPWR.n2 46.2505
R194 VPWR.n3 VPWR.n1 46.2505
R195 VPWR.n6 VPWR.n3 46.2505
R196 VPWR.n9 VPWR.n8 39.1534
R197 VPWR.n22 VPWR.n13 30.8711
R198 VPWR.n28 VPWR.n26 18.5005
R199 VPWR.n27 VPWR.n25 18.5005
R200 VPWR.n15 VPWR.n13 18.5005
R201 VPWR.n16 VPWR.n14 18.5005
R202 VPWR.n5 VPWR.n4 18.5005
R203 VPWR.n8 VPWR.n7 18.5005
R204 VPWR.n35 VPWR.n34 18.2416
R205 VPWR.n33 VPWR.n32 15.4172
R206 VPWR.n32 VPWR.n31 15.4172
R207 VPWR.n30 VPWR.n29 15.4172
R208 VPWR.n31 VPWR.n30 15.4172
R209 VPWR.n12 VPWR.n11 14.9974
R210 VPWR.n23 VPWR.t13 13.0025
R211 VPWR.n23 VPWR.t15 13.0025
R212 VPWR.n10 VPWR.t10 13.0025
R213 VPWR.n10 VPWR.t6 13.0025
R214 VPWR.n11 VPWR.n9 9.84217
R215 VPWR.n24 VPWR.n22 9.738
R216 VPWR.n35 VPWR.n24 9.39032
R217 VPWR.n12 VPWR 0.345167
R218 VPWR.n36 VPWR.n12 0.312267
R219 VPWR VPWR.n36 0.196333
R220 VPWR.n36 VPWR.n35 0.0459667
R221 ctrl.n0 ctrl.t1 649.289
R222 ctrl.n0 ctrl.t0 637.092
R223 ctrl.n1 ctrl.t2 312.086
R224 ctrl ctrl.n1 6.12074
R225 ctrl.n1 ctrl.n0 3.67146
C0 mod bus 5.87185f
C1 mod tgon_n 0.663384f
C2 bus tgon_n 0.929293f
C3 mod VPWR 1.14475f
C4 mod ctrl 0.030924f
C5 bus VPWR 0.879695f
C6 ctrl bus 0.090754f
C7 tgon_n VPWR 3.97533f
C8 ctrl tgon_n 0.699519f
C9 ctrl VPWR 0.903877f
C10 mod a_726_1810# 0.53907f
C11 bus a_726_1810# 0.207555f
C12 a_726_1810# tgon_n 0.565753f
C13 a_726_1810# VPWR 1.98842f
C14 ctrl a_726_1810# 0.002341f
C15 mod VGND 2.484136f
C16 bus VGND 1.194421f
C17 ctrl VGND 1.78843f
C18 VPWR VGND 11.995465f
C19 a_726_1810# VGND 2.64514f
C20 tgon_n VGND 5.100999f
C21 VPWR.n0 VGND 0.016773f
C22 VPWR.n1 VGND 0.018538f
C23 VPWR.n2 VGND 0.018538f
C24 VPWR.n3 VGND 0.018538f
C25 VPWR.n4 VGND 0.018228f
C26 VPWR.n5 VGND 0.115791f
C27 VPWR.t5 VGND 0.096069f
C28 VPWR.n6 VGND 0.038888f
C29 VPWR.t9 VGND 0.096069f
C30 VPWR.n7 VGND 0.115791f
C31 VPWR.n8 VGND 0.010682f
C32 VPWR.n9 VGND 0.010386f
C33 VPWR.t10 VGND 0.007126f
C34 VPWR.t6 VGND 0.007126f
C35 VPWR.n10 VGND 0.01887f
C36 VPWR.n11 VGND 0.165028f
C37 VPWR.n12 VGND 0.37261f
C38 VPWR.n13 VGND 0.01037f
C39 VPWR.n14 VGND 0.018228f
C40 VPWR.n15 VGND 0.115791f
C41 VPWR.n16 VGND 0.115791f
C42 VPWR.t12 VGND 0.096069f
C43 VPWR.t14 VGND 0.096069f
C44 VPWR.n17 VGND 0.018538f
C45 VPWR.n18 VGND 0.018538f
C46 VPWR.n19 VGND 0.038888f
C47 VPWR.n20 VGND 0.018538f
C48 VPWR.n21 VGND 0.017105f
C49 VPWR.n22 VGND 0.010215f
C50 VPWR.t13 VGND 0.007126f
C51 VPWR.t15 VGND 0.007126f
C52 VPWR.n23 VGND 0.015796f
C53 VPWR.n24 VGND 0.060276f
C54 VPWR.n25 VGND 0.02366f
C55 VPWR.n26 VGND 0.026896f
C56 VPWR.n27 VGND 0.124459f
C57 VPWR.n28 VGND 0.124459f
C58 VPWR.t2 VGND 0.115513f
C59 VPWR.t11 VGND 0.077776f
C60 VPWR.t7 VGND 0.077776f
C61 VPWR.t3 VGND 0.058332f
C62 VPWR.n29 VGND 0.026786f
C63 VPWR.n30 VGND 0.026786f
C64 VPWR.t1 VGND 0.115513f
C65 VPWR.t4 VGND 0.077776f
C66 VPWR.t8 VGND 0.077776f
C67 VPWR.t0 VGND 0.058332f
C68 VPWR.n31 VGND 0.038888f
C69 VPWR.n32 VGND 0.026786f
C70 VPWR.n33 VGND 0.01638f
C71 VPWR.n34 VGND 0.025372f
C72 VPWR.n35 VGND 0.5165f
C73 VPWR.n36 VGND 0.268652f
C74 tgon_n.n0 VGND 0.13977f
C75 tgon_n.n1 VGND 0.292124f
C76 tgon_n.n2 VGND 0.13887f
C77 tgon_n.n3 VGND 0.227825f
C78 tgon_n.t5 VGND 0.05008f
C79 tgon_n.t8 VGND 0.057588f
C80 tgon_n.n4 VGND 0.698154f
C81 tgon_n.t4 VGND 0.053894f
C82 tgon_n.t11 VGND 0.050065f
C83 tgon_n.t7 VGND 0.050024f
C84 tgon_n.t13 VGND 0.050024f
C85 tgon_n.t9 VGND 0.050024f
C86 tgon_n.t3 VGND 0.050064f
C87 tgon_n.t10 VGND 0.050024f
C88 tgon_n.t6 VGND 0.050024f
C89 tgon_n.t12 VGND 0.050039f
C90 tgon_n.n5 VGND 0.354803f
C91 tgon_n.t1 VGND 0.112162f
C92 tgon_n.t2 VGND 0.111578f
C93 tgon_n.n6 VGND 0.341162f
C94 tgon_n.t0 VGND 0.094881f
C95 bus.t3 VGND 0.23176f
C96 bus.t0 VGND 0.063362f
C97 bus.t4 VGND 0.063362f
C98 bus.n0 VGND 0.143272f
C99 bus.n1 VGND 0.709642f
C100 bus.t1 VGND 0.063362f
C101 bus.t5 VGND 0.063362f
C102 bus.n2 VGND 0.143444f
C103 bus.n3 VGND 0.358564f
C104 bus.t11 VGND 0.063362f
C105 bus.t6 VGND 0.063362f
C106 bus.n4 VGND 0.143444f
C107 bus.n5 VGND 0.357489f
C108 bus.t2 VGND 0.230512f
C109 bus.n6 VGND 0.697744f
C110 bus.t7 VGND 0.063362f
C111 bus.t10 VGND 0.063362f
C112 bus.n7 VGND 0.134142f
C113 bus.t9 VGND 0.063362f
C114 bus.t8 VGND 0.063362f
C115 bus.n8 VGND 0.13294f
C116 bus.n9 VGND 0.281674f
C117 bus.n10 VGND 0.562805f
C118 bus.n11 VGND 0.862466f
C119 mod.t8 VGND 0.180421f
C120 mod.t10 VGND 0.047388f
C121 mod.t7 VGND 0.047388f
C122 mod.n0 VGND 0.12683f
C123 mod.n1 VGND 0.53618f
C124 mod.t9 VGND 0.178441f
C125 mod.n2 VGND 0.541748f
C126 mod.t6 VGND 0.047388f
C127 mod.t2 VGND 0.047388f
C128 mod.n3 VGND 0.104848f
C129 mod.t5 VGND 0.047388f
C130 mod.t11 VGND 0.047388f
C131 mod.n4 VGND 0.103964f
C132 mod.n5 VGND 0.479416f
C133 mod.t4 VGND 0.047388f
C134 mod.t1 VGND 0.047388f
C135 mod.n6 VGND 0.104027f
C136 mod.n7 VGND 0.230276f
C137 mod.t3 VGND 0.047388f
C138 mod.t0 VGND 0.047388f
C139 mod.n8 VGND 0.104154f
C140 mod.n9 VGND 0.297699f
C141 mod.n10 VGND 1.36749f
C142 mod.n11 VGND 0.863838f
.ends

