magic
tech sky130A
magscale 1 2
timestamp 1712309281
<< nwell >>
rect -720 -519 720 519
<< pmoslvt >>
rect -524 -300 -424 300
rect -366 -300 -266 300
rect -208 -300 -108 300
rect -50 -300 50 300
rect 108 -300 208 300
rect 266 -300 366 300
rect 424 -300 524 300
<< pdiff >>
rect -582 288 -524 300
rect -582 -288 -570 288
rect -536 -288 -524 288
rect -582 -300 -524 -288
rect -424 288 -366 300
rect -424 -288 -412 288
rect -378 -288 -366 288
rect -424 -300 -366 -288
rect -266 288 -208 300
rect -266 -288 -254 288
rect -220 -288 -208 288
rect -266 -300 -208 -288
rect -108 288 -50 300
rect -108 -288 -96 288
rect -62 -288 -50 288
rect -108 -300 -50 -288
rect 50 288 108 300
rect 50 -288 62 288
rect 96 -288 108 288
rect 50 -300 108 -288
rect 208 288 266 300
rect 208 -288 220 288
rect 254 -288 266 288
rect 208 -300 266 -288
rect 366 288 424 300
rect 366 -288 378 288
rect 412 -288 424 288
rect 366 -300 424 -288
rect 524 288 582 300
rect 524 -288 536 288
rect 570 -288 582 288
rect 524 -300 582 -288
<< pdiffc >>
rect -570 -288 -536 288
rect -412 -288 -378 288
rect -254 -288 -220 288
rect -96 -288 -62 288
rect 62 -288 96 288
rect 220 -288 254 288
rect 378 -288 412 288
rect 536 -288 570 288
<< nsubdiff >>
rect -684 449 -588 483
rect 588 449 684 483
rect -684 387 -650 449
rect 650 387 684 449
rect -684 -449 -650 -387
rect 650 -449 684 -387
rect -684 -483 -588 -449
rect 588 -483 684 -449
<< nsubdiffcont >>
rect -588 449 588 483
rect -684 -387 -650 387
rect 650 -387 684 387
rect -588 -483 588 -449
<< poly >>
rect -524 381 -424 397
rect -524 347 -508 381
rect -440 347 -424 381
rect -524 300 -424 347
rect -366 381 -266 397
rect -366 347 -350 381
rect -282 347 -266 381
rect -366 300 -266 347
rect -208 381 -108 397
rect -208 347 -192 381
rect -124 347 -108 381
rect -208 300 -108 347
rect -50 381 50 397
rect -50 347 -34 381
rect 34 347 50 381
rect -50 300 50 347
rect 108 381 208 397
rect 108 347 124 381
rect 192 347 208 381
rect 108 300 208 347
rect 266 381 366 397
rect 266 347 282 381
rect 350 347 366 381
rect 266 300 366 347
rect 424 381 524 397
rect 424 347 440 381
rect 508 347 524 381
rect 424 300 524 347
rect -524 -347 -424 -300
rect -524 -381 -508 -347
rect -440 -381 -424 -347
rect -524 -397 -424 -381
rect -366 -347 -266 -300
rect -366 -381 -350 -347
rect -282 -381 -266 -347
rect -366 -397 -266 -381
rect -208 -347 -108 -300
rect -208 -381 -192 -347
rect -124 -381 -108 -347
rect -208 -397 -108 -381
rect -50 -347 50 -300
rect -50 -381 -34 -347
rect 34 -381 50 -347
rect -50 -397 50 -381
rect 108 -347 208 -300
rect 108 -381 124 -347
rect 192 -381 208 -347
rect 108 -397 208 -381
rect 266 -347 366 -300
rect 266 -381 282 -347
rect 350 -381 366 -347
rect 266 -397 366 -381
rect 424 -347 524 -300
rect 424 -381 440 -347
rect 508 -381 524 -347
rect 424 -397 524 -381
<< polycont >>
rect -508 347 -440 381
rect -350 347 -282 381
rect -192 347 -124 381
rect -34 347 34 381
rect 124 347 192 381
rect 282 347 350 381
rect 440 347 508 381
rect -508 -381 -440 -347
rect -350 -381 -282 -347
rect -192 -381 -124 -347
rect -34 -381 34 -347
rect 124 -381 192 -347
rect 282 -381 350 -347
rect 440 -381 508 -347
<< locali >>
rect -684 449 -588 483
rect 588 449 684 483
rect -684 387 -650 449
rect 650 387 684 449
rect -524 347 -508 381
rect -440 347 -424 381
rect -366 347 -350 381
rect -282 347 -266 381
rect -208 347 -192 381
rect -124 347 -108 381
rect -50 347 -34 381
rect 34 347 50 381
rect 108 347 124 381
rect 192 347 208 381
rect 266 347 282 381
rect 350 347 366 381
rect 424 347 440 381
rect 508 347 524 381
rect -570 288 -536 304
rect -570 -304 -536 -288
rect -412 288 -378 304
rect -412 -304 -378 -288
rect -254 288 -220 304
rect -254 -304 -220 -288
rect -96 288 -62 304
rect -96 -304 -62 -288
rect 62 288 96 304
rect 62 -304 96 -288
rect 220 288 254 304
rect 220 -304 254 -288
rect 378 288 412 304
rect 378 -304 412 -288
rect 536 288 570 304
rect 536 -304 570 -288
rect -524 -381 -508 -347
rect -440 -381 -424 -347
rect -366 -381 -350 -347
rect -282 -381 -266 -347
rect -208 -381 -192 -347
rect -124 -381 -108 -347
rect -50 -381 -34 -347
rect 34 -381 50 -347
rect 108 -381 124 -347
rect 192 -381 208 -347
rect 266 -381 282 -347
rect 350 -381 366 -347
rect 424 -381 440 -347
rect 508 -381 524 -347
rect -684 -449 -650 -387
rect 650 -449 684 -387
rect -684 -483 -588 -449
rect 588 -483 684 -449
<< viali >>
rect -508 347 -440 381
rect -350 347 -282 381
rect -192 347 -124 381
rect -34 347 34 381
rect 124 347 192 381
rect 282 347 350 381
rect 440 347 508 381
rect -570 -288 -536 288
rect -412 -288 -378 288
rect -254 -288 -220 288
rect -96 -288 -62 288
rect 62 -288 96 288
rect 220 -288 254 288
rect 378 -288 412 288
rect 536 -288 570 288
rect -508 -381 -440 -347
rect -350 -381 -282 -347
rect -192 -381 -124 -347
rect -34 -381 34 -347
rect 124 -381 192 -347
rect 282 -381 350 -347
rect 440 -381 508 -347
<< metal1 >>
rect -520 381 -428 387
rect -520 347 -508 381
rect -440 347 -428 381
rect -520 341 -428 347
rect -362 381 -270 387
rect -362 347 -350 381
rect -282 347 -270 381
rect -362 341 -270 347
rect -204 381 -112 387
rect -204 347 -192 381
rect -124 347 -112 381
rect -204 341 -112 347
rect -46 381 46 387
rect -46 347 -34 381
rect 34 347 46 381
rect -46 341 46 347
rect 112 381 204 387
rect 112 347 124 381
rect 192 347 204 381
rect 112 341 204 347
rect 270 381 362 387
rect 270 347 282 381
rect 350 347 362 381
rect 270 341 362 347
rect 428 381 520 387
rect 428 347 440 381
rect 508 347 520 381
rect 428 341 520 347
rect -576 288 -530 300
rect -576 -288 -570 288
rect -536 -288 -530 288
rect -576 -300 -530 -288
rect -418 288 -372 300
rect -418 -288 -412 288
rect -378 -288 -372 288
rect -418 -300 -372 -288
rect -260 288 -214 300
rect -260 -288 -254 288
rect -220 -288 -214 288
rect -260 -300 -214 -288
rect -102 288 -56 300
rect -102 -288 -96 288
rect -62 -288 -56 288
rect -102 -300 -56 -288
rect 56 288 102 300
rect 56 -288 62 288
rect 96 -288 102 288
rect 56 -300 102 -288
rect 214 288 260 300
rect 214 -288 220 288
rect 254 -288 260 288
rect 214 -300 260 -288
rect 372 288 418 300
rect 372 -288 378 288
rect 412 -288 418 288
rect 372 -300 418 -288
rect 530 288 576 300
rect 530 -288 536 288
rect 570 -288 576 288
rect 530 -300 576 -288
rect -520 -347 -428 -341
rect -520 -381 -508 -347
rect -440 -381 -428 -347
rect -520 -387 -428 -381
rect -362 -347 -270 -341
rect -362 -381 -350 -347
rect -282 -381 -270 -347
rect -362 -387 -270 -381
rect -204 -347 -112 -341
rect -204 -381 -192 -347
rect -124 -381 -112 -347
rect -204 -387 -112 -381
rect -46 -347 46 -341
rect -46 -381 -34 -347
rect 34 -381 46 -347
rect -46 -387 46 -381
rect 112 -347 204 -341
rect 112 -381 124 -347
rect 192 -381 204 -347
rect 112 -387 204 -381
rect 270 -347 362 -341
rect 270 -381 282 -347
rect 350 -381 362 -347
rect 270 -387 362 -381
rect 428 -347 520 -341
rect 428 -381 440 -347
rect 508 -381 520 -347
rect 428 -387 520 -381
<< properties >>
string FIXED_BBOX -667 -466 667 466
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 3 l 0.5 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
