magic
tech sky130A
magscale 1 2
timestamp 1711023331
<< error_s >>
rect 2382 3882 2440 3888
rect 2574 3882 2632 3888
rect 2382 3848 2394 3882
rect 2574 3848 2586 3882
rect 2382 3842 2440 3848
rect 2574 3842 2632 3848
rect 2286 3272 2344 3278
rect 2478 3272 2536 3278
rect 2286 3238 2298 3272
rect 2478 3238 2490 3272
rect 2286 3232 2344 3238
rect 2478 3232 2536 3238
rect 682 3172 740 3178
rect 1286 3172 1344 3178
rect 682 3138 694 3172
rect 1286 3138 1298 3172
rect 682 3132 740 3138
rect 1286 3132 1344 3138
rect 2382 2800 2440 2806
rect 2574 2800 2632 2806
rect 2766 2800 2824 2806
rect 2958 2800 3016 2806
rect 2382 2766 2394 2800
rect 2574 2766 2586 2800
rect 2766 2766 2778 2800
rect 2958 2766 2970 2800
rect 2382 2760 2440 2766
rect 2574 2760 2632 2766
rect 2766 2760 2824 2766
rect 2958 2760 3016 2766
rect 1382 2400 1440 2406
rect 682 2382 740 2388
rect 682 2348 694 2382
rect 1382 2366 1394 2400
rect 1382 2360 1440 2366
rect 682 2342 740 2348
rect 2286 2172 2344 2178
rect 2478 2172 2536 2178
rect 2670 2172 2728 2178
rect 2862 2172 2920 2178
rect 2286 2138 2298 2172
rect 2478 2138 2490 2172
rect 2670 2138 2682 2172
rect 2862 2138 2874 2172
rect 2286 2132 2344 2138
rect 2478 2132 2536 2138
rect 2670 2132 2728 2138
rect 2862 2132 2920 2138
rect 682 1772 740 1778
rect 1286 1772 1344 1778
rect 682 1738 694 1772
rect 1286 1738 1298 1772
rect 682 1732 740 1738
rect 1286 1732 1344 1738
<< pwell >>
rect 970 3450 1060 3510
<< metal1 >>
rect 684 3970 690 4030
rect 750 3970 756 4030
rect 690 3910 1440 3970
rect 690 3740 750 3910
rect 1380 3750 1440 3910
rect 415 3451 421 3510
rect 480 3451 689 3510
rect 730 3450 1290 3510
rect 1430 3450 1780 3510
rect 1840 3450 1846 3510
<< via1 >>
rect 690 3970 750 4030
rect 421 3451 480 3510
rect 1780 3450 1840 3510
<< metal2 >>
rect 690 4108 750 4110
rect 683 4052 692 4108
rect 748 4052 757 4108
rect 690 4030 750 4052
rect 690 3964 750 3970
rect 272 3451 281 3511
rect 341 3510 350 3511
rect 421 3510 480 3516
rect 341 3451 421 3510
rect 421 3445 480 3451
rect 1780 3510 1840 3516
rect 1840 3450 1880 3510
rect 1940 3450 1949 3510
rect 1780 3444 1840 3450
<< via2 >>
rect 692 4052 748 4108
rect 281 3451 341 3511
rect 1880 3450 1940 3510
<< metal3 >>
rect 120 4346 360 4352
rect 120 2358 126 4346
rect 354 2358 360 4346
rect 687 4110 753 4113
rect 890 4110 950 4352
rect 687 4108 950 4110
rect 687 4052 692 4108
rect 748 4052 950 4108
rect 687 4050 950 4052
rect 1750 4346 1930 4352
rect 687 4047 753 4050
rect 1750 3958 1756 4346
rect 1924 3958 1930 4346
rect 1750 3952 1930 3958
rect 3320 4346 3560 4352
rect 1875 3510 1945 3515
rect 3320 3510 3326 4346
rect 1875 3450 1880 3510
rect 1940 3450 3326 3510
rect 1875 3445 1945 3450
rect 120 2352 360 2358
rect 1750 2746 1930 2752
rect 1750 2358 1756 2746
rect 1924 2358 1930 2746
rect 1750 2352 1930 2358
rect 3320 2358 3326 3450
rect 3554 2358 3560 4346
rect 3320 2352 3560 2358
<< via3 >>
rect 126 3511 354 4346
rect 126 3451 281 3511
rect 281 3451 341 3511
rect 341 3451 354 3511
rect 126 2358 354 3451
rect 1756 3958 1924 4346
rect 1756 2358 1924 2746
rect 3326 2358 3554 4346
<< metal4 >>
rect 120 4346 360 4352
rect 120 2358 126 4346
rect 354 2358 360 4346
rect 1750 4346 1930 4352
rect 1750 3958 1756 4346
rect 1924 3958 1930 4346
rect 1750 3952 1930 3958
rect 3320 4346 3560 4352
rect 120 0 360 2358
rect 1750 2746 1930 2752
rect 1750 2358 1756 2746
rect 1924 2358 1930 2746
rect 1750 2352 1930 2358
rect 3320 2358 3326 4346
rect 3554 2358 3560 4346
rect 3320 0 3560 2358
use sky130_fd_pr__nfet_01v8_H7HSAV  XM1
timestamp 1711022820
transform 1 0 711 0 1 3460
box -211 -460 211 460
use sky130_fd_pr__pfet_01v8_XJT9DL  XM2
timestamp 1711022820
transform 1 0 1363 0 1 3469
box -263 -469 263 469
use sky130_fd_pr__nfet_01v8_5ZNSAF  XM3
timestamp 1711022820
transform 1 0 2459 0 1 3560
box -359 -460 359 460
use sky130_fd_pr__pfet_01v8_XJKGNP  XM4A
timestamp 1711022820
transform 1 0 2651 0 1 2469
box -551 -469 551 469
use sky130_fd_pr__pfet_01v8_XJT9DL  XM4
timestamp 1711022820
transform 1 0 1363 0 1 2069
box -263 -469 263 469
use sky130_fd_pr__nfet_01v8_H7HSAV  XM5
timestamp 1711022820
transform 1 0 711 0 1 2060
box -211 -460 211 460
<< labels >>
rlabel metal4 3320 0 3560 4352 1 VPWR
port 2 n power input
rlabel metal4 1750 3952 1930 4352 1 mod
port 3 n analog bidirectional
rlabel metal4 1750 2352 1930 2752 1 bus
port 4 n analog bidirectional
rlabel metal3 890 4172 950 4352 1 ctrl
port 5 n signal input
rlabel metal4 120 0 360 4352 1 VGND
port 1 n ground input
<< properties >>
string FIXED_BBOX 0 0 3680 4352
<< end >>
