VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_asw_1v8
  CLASS BLOCK ;
  FOREIGN tt_asw_1v8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.400 BY 21.760 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.600 0.000 1.800 21.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.600 0.000 17.800 21.760 ;
    END
  END VPWR
  PIN mod
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 8.750 19.760 9.650 21.760 ;
    END
  END mod
  PIN bus
    DIRECTION INOUT ;
    USE ANALOG ;
    PORT
      LAYER met4 ;
        RECT 8.750 11.760 9.650 13.760 ;
    END
  END bus
  PIN ctrl
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4.450 20.860 4.750 21.760 ;
    END
  END ctrl
  OBS
      LAYER pwell ;
        RECT 3.190 2.720 5.650 14.820 ;
      LAYER nwell ;
        RECT 6.210 10.540 8.670 22.730 ;
        RECT 12.880 10.470 15.340 22.660 ;
      LAYER pwell ;
        RECT 6.570 6.660 9.030 9.760 ;
      LAYER nwell ;
        RECT 6.890 1.270 9.350 5.460 ;
      LAYER pwell ;
        RECT 10.380 1.580 12.840 4.680 ;
      LAYER nwell ;
        RECT 12.905 1.145 15.365 5.335 ;
      LAYER li1 ;
        RECT 6.390 22.380 8.490 22.550 ;
        RECT 3.370 14.470 5.470 14.640 ;
        RECT 3.370 3.070 3.540 14.470 ;
        RECT 4.170 13.960 4.670 14.130 ;
        RECT 3.940 3.750 4.110 13.790 ;
        RECT 4.730 3.750 4.900 13.790 ;
        RECT 4.170 3.410 4.670 3.580 ;
        RECT 5.300 3.070 5.470 14.470 ;
        RECT 6.390 10.890 6.560 22.380 ;
        RECT 7.190 21.870 7.690 22.040 ;
        RECT 6.960 11.615 7.130 21.655 ;
        RECT 7.750 11.615 7.920 21.655 ;
        RECT 7.190 11.230 7.690 11.400 ;
        RECT 8.320 10.890 8.490 22.380 ;
        RECT 6.390 10.720 8.490 10.890 ;
        RECT 13.060 22.310 15.160 22.480 ;
        RECT 13.060 10.820 13.230 22.310 ;
        RECT 13.860 21.800 14.360 21.970 ;
        RECT 13.630 11.545 13.800 21.585 ;
        RECT 14.420 11.545 14.590 21.585 ;
        RECT 13.860 11.160 14.360 11.330 ;
        RECT 14.990 10.820 15.160 22.310 ;
        RECT 13.060 10.650 15.160 10.820 ;
        RECT 6.750 9.410 8.850 9.580 ;
        RECT 6.750 7.010 6.920 9.410 ;
        RECT 7.550 8.900 8.050 9.070 ;
        RECT 7.320 7.690 7.490 8.730 ;
        RECT 8.110 7.690 8.280 8.730 ;
        RECT 7.550 7.350 8.050 7.520 ;
        RECT 8.680 7.010 8.850 9.410 ;
        RECT 6.750 6.840 8.850 7.010 ;
        RECT 3.370 2.900 5.470 3.070 ;
        RECT 7.070 5.110 9.170 5.280 ;
        RECT 7.070 1.620 7.240 5.110 ;
        RECT 7.870 4.600 8.370 4.770 ;
        RECT 7.640 2.345 7.810 4.385 ;
        RECT 8.430 2.345 8.600 4.385 ;
        RECT 7.870 1.960 8.370 2.130 ;
        RECT 9.000 1.620 9.170 5.110 ;
        RECT 13.085 4.985 15.185 5.155 ;
        RECT 10.560 4.330 12.660 4.500 ;
        RECT 10.560 1.930 10.730 4.330 ;
        RECT 11.360 3.820 11.860 3.990 ;
        RECT 11.130 2.610 11.300 3.650 ;
        RECT 11.920 2.610 12.090 3.650 ;
        RECT 11.360 2.270 11.860 2.440 ;
        RECT 12.490 1.930 12.660 4.330 ;
        RECT 10.560 1.760 12.660 1.930 ;
        RECT 7.070 1.450 9.170 1.620 ;
        RECT 13.085 1.495 13.255 4.985 ;
        RECT 13.885 4.475 14.385 4.645 ;
        RECT 13.655 2.220 13.825 4.260 ;
        RECT 14.445 2.220 14.615 4.260 ;
        RECT 13.885 1.835 14.385 2.005 ;
        RECT 15.015 1.495 15.185 4.985 ;
        RECT 13.085 1.325 15.185 1.495 ;
      LAYER mcon ;
        RECT 4.250 13.960 4.590 14.130 ;
        RECT 3.940 3.830 4.110 13.710 ;
        RECT 4.730 3.830 4.900 13.710 ;
        RECT 4.250 3.410 4.590 3.580 ;
        RECT 7.270 21.870 7.610 22.040 ;
        RECT 6.960 11.695 7.130 21.575 ;
        RECT 7.750 11.695 7.920 21.575 ;
        RECT 7.270 11.230 7.610 11.400 ;
        RECT 13.940 21.800 14.280 21.970 ;
        RECT 13.630 11.625 13.800 21.505 ;
        RECT 14.420 11.625 14.590 21.505 ;
        RECT 13.940 11.160 14.280 11.330 ;
        RECT 7.630 8.900 7.970 9.070 ;
        RECT 7.320 7.770 7.490 8.650 ;
        RECT 8.110 7.770 8.280 8.650 ;
        RECT 7.630 7.350 7.970 7.520 ;
        RECT 7.950 4.600 8.290 4.770 ;
        RECT 7.640 2.425 7.810 4.305 ;
        RECT 8.430 2.425 8.600 4.305 ;
        RECT 7.950 1.960 8.290 2.130 ;
        RECT 11.440 3.820 11.780 3.990 ;
        RECT 11.130 2.690 11.300 3.570 ;
        RECT 11.920 2.690 12.090 3.570 ;
        RECT 11.440 2.270 11.780 2.440 ;
        RECT 13.965 4.475 14.305 4.645 ;
        RECT 13.655 2.300 13.825 4.180 ;
        RECT 14.445 2.300 14.615 4.180 ;
        RECT 13.965 1.835 14.305 2.005 ;
      LAYER met1 ;
        RECT 7.210 21.840 7.670 22.070 ;
        RECT 13.880 21.770 14.340 22.000 ;
        RECT 4.190 13.930 4.650 14.160 ;
        RECT 3.910 3.770 4.140 13.770 ;
        RECT 4.700 3.770 4.930 13.770 ;
        RECT 6.930 11.635 7.160 21.635 ;
        RECT 7.720 11.635 7.950 21.635 ;
        RECT 13.600 11.565 13.830 21.565 ;
        RECT 14.390 11.565 14.620 21.565 ;
        RECT 7.210 11.200 7.670 11.430 ;
        RECT 13.880 11.130 14.340 11.360 ;
        RECT 7.570 8.870 8.030 9.100 ;
        RECT 7.290 7.710 7.520 8.710 ;
        RECT 8.080 7.710 8.310 8.710 ;
        RECT 7.570 7.320 8.030 7.550 ;
        RECT 7.890 4.570 8.350 4.800 ;
        RECT 13.905 4.445 14.365 4.675 ;
        RECT 4.190 3.380 4.650 3.610 ;
        RECT 7.610 2.365 7.840 4.365 ;
        RECT 8.400 2.365 8.630 4.365 ;
        RECT 11.380 3.790 11.840 4.020 ;
        RECT 11.100 2.630 11.330 3.630 ;
        RECT 11.890 2.630 12.120 3.630 ;
        RECT 11.380 2.240 11.840 2.470 ;
        RECT 13.625 2.240 13.855 4.240 ;
        RECT 14.415 2.240 14.645 4.240 ;
        RECT 7.890 1.930 8.350 2.160 ;
        RECT 13.905 1.805 14.365 2.035 ;
      LAYER met3 ;
        RECT 0.600 11.760 1.800 21.760 ;
        RECT 8.750 19.760 9.650 21.760 ;
        RECT 8.750 11.760 9.650 13.760 ;
        RECT 16.600 11.760 17.800 21.760 ;
      LAYER via3 ;
        RECT 0.630 11.790 1.770 21.730 ;
        RECT 8.780 19.790 9.620 21.730 ;
        RECT 8.780 11.790 9.620 13.730 ;
        RECT 16.630 11.790 17.770 21.730 ;
  END
END tt_asw_1v8
END LIBRARY

