magic
tech sky130A
magscale 1 2
timestamp 1712328979
<< locali >>
rect 120 4332 3560 4352
rect 120 4132 140 4332
rect 340 4156 3560 4332
rect 340 4132 400 4156
rect 120 4122 400 4132
rect 3540 4122 3560 4156
rect 120 4020 3560 4122
rect 1016 3790 1910 4020
rect 1996 2664 3364 2900
rect 120 2582 3560 2664
rect 120 2548 140 2582
rect 3280 2572 3560 2582
rect 3280 2548 3340 2572
rect 120 2372 3340 2548
rect 3540 2372 3560 2572
rect 120 2352 3560 2372
<< viali >>
rect 140 4132 340 4332
rect 400 4122 3540 4156
rect 604 3594 638 3870
rect 692 3594 726 3870
rect 604 2825 638 3101
rect 700 2825 734 3101
rect 796 2825 830 3101
rect 140 2548 3280 2582
rect 3340 2372 3540 2572
<< metal1 >>
rect 120 4332 3560 4352
rect 120 4132 140 4332
rect 340 4156 598 4332
rect 650 4156 3560 4332
rect 340 4132 400 4156
rect 120 4122 400 4132
rect 3540 4122 3560 4156
rect 120 4112 3560 4122
rect 190 3912 378 3962
rect 506 3912 694 3962
rect 190 3552 236 3912
rect 282 3876 334 3882
rect 282 3582 334 3588
rect 364 3876 416 3882
rect 364 3582 416 3588
rect 506 3552 552 3912
rect 598 3876 650 3882
rect 598 3582 650 3588
rect 680 3876 732 3882
rect 680 3582 732 3588
rect 1028 3682 1746 3728
rect 2008 3690 3204 3736
rect 190 3502 378 3552
rect 506 3502 694 3552
rect 190 3388 236 3502
rect 184 3382 242 3388
rect 506 3384 552 3502
rect 1028 3384 1074 3682
rect 1120 3642 1174 3650
rect 184 3316 242 3322
rect 502 3378 556 3384
rect 1024 3378 1078 3384
rect 556 3332 940 3372
rect 502 3320 556 3326
rect 190 3202 236 3316
rect 506 3202 552 3320
rect 86 3152 380 3202
rect 506 3152 800 3202
rect 86 2774 132 3152
rect 178 3108 230 3114
rect 178 2812 230 2818
rect 270 3108 324 3114
rect 270 2812 324 2818
rect 364 3108 416 3114
rect 364 2812 416 2818
rect 506 2774 552 3152
rect 598 3108 650 3114
rect 598 2812 650 2818
rect 690 3108 744 3114
rect 690 2812 744 2818
rect 784 3108 836 3114
rect 900 2920 940 3332
rect 1024 3320 1078 3326
rect 1028 3018 1074 3320
rect 1120 3048 1174 3056
rect 1278 3642 1332 3650
rect 1278 3048 1332 3056
rect 1436 3642 1490 3650
rect 1436 3048 1490 3056
rect 1594 3642 1648 3650
rect 1594 3048 1648 3056
rect 1752 3642 1806 3650
rect 2008 3372 2054 3690
rect 1752 3048 1806 3056
rect 1900 3332 2054 3372
rect 1028 2972 1746 3018
rect 1900 2920 1940 3332
rect 2008 3008 2054 3332
rect 2100 3642 2154 3650
rect 2100 3048 2154 3056
rect 2258 3642 2312 3650
rect 2258 3048 2312 3056
rect 2416 3642 2470 3650
rect 2416 3048 2470 3056
rect 2574 3642 2628 3650
rect 2574 3048 2628 3056
rect 2732 3642 2786 3650
rect 2732 3048 2786 3056
rect 2890 3642 2944 3650
rect 2890 3048 2944 3056
rect 3048 3642 3102 3650
rect 3048 3048 3102 3056
rect 3206 3642 3260 3650
rect 3206 3048 3260 3056
rect 2008 2962 3204 3008
rect 900 2880 1940 2920
rect 784 2812 836 2818
rect 86 2724 380 2774
rect 506 2724 800 2774
rect 120 2582 3560 2592
rect 120 2548 140 2582
rect 3280 2572 3560 2582
rect 3280 2548 3340 2572
rect 120 2372 178 2548
rect 230 2372 364 2548
rect 416 2372 598 2548
rect 650 2372 784 2548
rect 836 2372 3340 2548
rect 3540 2372 3560 2572
rect 120 2352 3560 2372
<< via1 >>
rect 140 4132 340 4332
rect 598 4156 650 4332
rect 598 4132 650 4156
rect 282 3588 334 3876
rect 364 3588 416 3876
rect 598 3870 650 3876
rect 598 3594 604 3870
rect 604 3594 638 3870
rect 638 3594 650 3870
rect 598 3588 650 3594
rect 680 3870 732 3876
rect 680 3594 692 3870
rect 692 3594 726 3870
rect 726 3594 732 3870
rect 680 3588 732 3594
rect 184 3322 242 3382
rect 502 3326 556 3378
rect 178 2818 230 3108
rect 270 2818 324 3108
rect 364 2818 416 3108
rect 598 3101 650 3108
rect 598 2825 604 3101
rect 604 2825 638 3101
rect 638 2825 650 3101
rect 598 2818 650 2825
rect 690 3101 744 3108
rect 690 2825 700 3101
rect 700 2825 734 3101
rect 734 2825 744 3101
rect 690 2818 744 2825
rect 784 3101 836 3108
rect 784 2825 796 3101
rect 796 2825 830 3101
rect 830 2825 836 3101
rect 1024 3326 1078 3378
rect 1120 3056 1174 3642
rect 1278 3056 1332 3642
rect 1436 3056 1490 3642
rect 1594 3056 1648 3642
rect 1752 3056 1806 3642
rect 2100 3056 2154 3642
rect 2258 3056 2312 3642
rect 2416 3056 2470 3642
rect 2574 3056 2628 3642
rect 2732 3056 2786 3642
rect 2890 3056 2944 3642
rect 3048 3056 3102 3642
rect 3206 3056 3260 3642
rect 784 2818 836 2825
rect 178 2548 230 2572
rect 364 2548 416 2572
rect 598 2548 650 2572
rect 784 2548 836 2572
rect 178 2372 230 2548
rect 364 2372 416 2548
rect 598 2372 650 2548
rect 784 2372 836 2548
rect 3340 2372 3540 2572
<< metal2 >>
rect 120 4332 360 4352
rect 120 4132 140 4332
rect 340 4132 360 4332
rect 120 4112 360 4132
rect 598 4332 650 4352
rect 282 3876 334 4112
rect 282 3582 334 3588
rect 364 3876 416 3882
rect 184 3382 242 3392
rect 364 3372 416 3588
rect 598 3876 650 4132
rect 598 3582 650 3588
rect 680 3876 732 3882
rect 496 3372 502 3378
rect 184 3312 242 3322
rect 270 3332 502 3372
rect 178 3108 230 3114
rect 178 2572 230 2818
rect 270 3108 324 3332
rect 496 3326 502 3332
rect 556 3326 562 3378
rect 680 3372 732 3588
rect 1118 3642 1176 3652
rect 1018 3372 1024 3378
rect 680 3332 1024 3372
rect 270 2812 324 2818
rect 364 3108 416 3114
rect 178 2352 230 2372
rect 364 2572 416 2818
rect 364 2352 416 2372
rect 598 3108 650 3114
rect 598 2572 650 2818
rect 690 3108 744 3332
rect 1018 3326 1024 3332
rect 1078 3326 1084 3378
rect 690 2812 744 2818
rect 784 3108 836 3114
rect 1118 3046 1176 3056
rect 1276 3642 1334 3652
rect 1276 3046 1334 3056
rect 1434 3642 1492 3652
rect 1434 3046 1492 3056
rect 1592 3642 1650 3652
rect 1592 3046 1650 3056
rect 1750 3642 1808 3652
rect 1750 3046 1808 3056
rect 2098 3642 2156 3652
rect 2098 3046 2156 3056
rect 2256 3642 2314 3652
rect 2256 3046 2314 3056
rect 2414 3642 2472 3652
rect 2414 3046 2472 3056
rect 2572 3642 2630 3652
rect 2572 3046 2630 3056
rect 2730 3642 2788 3652
rect 2730 3046 2788 3056
rect 2888 3642 2946 3652
rect 2888 3046 2946 3056
rect 3046 3642 3104 3652
rect 3046 3046 3104 3056
rect 3204 3642 3262 3652
rect 3204 3046 3262 3056
rect 598 2352 650 2372
rect 784 2572 836 2818
rect 784 2352 836 2372
rect 3320 2572 3560 2592
rect 3320 2372 3340 2572
rect 3540 2372 3560 2572
rect 3320 2352 3560 2372
<< via2 >>
rect 140 4132 340 4332
rect 184 3322 242 3382
rect 1118 3056 1120 3642
rect 1120 3056 1174 3642
rect 1174 3056 1176 3642
rect 1276 3056 1278 3642
rect 1278 3056 1332 3642
rect 1332 3056 1334 3642
rect 1434 3056 1436 3642
rect 1436 3056 1490 3642
rect 1490 3056 1492 3642
rect 1592 3056 1594 3642
rect 1594 3056 1648 3642
rect 1648 3056 1650 3642
rect 1750 3056 1752 3642
rect 1752 3056 1806 3642
rect 1806 3056 1808 3642
rect 2098 3056 2100 3642
rect 2100 3056 2154 3642
rect 2154 3056 2156 3642
rect 2256 3056 2258 3642
rect 2258 3056 2312 3642
rect 2312 3056 2314 3642
rect 2414 3056 2416 3642
rect 2416 3056 2470 3642
rect 2470 3056 2472 3642
rect 2572 3056 2574 3642
rect 2574 3056 2628 3642
rect 2628 3056 2630 3642
rect 2730 3056 2732 3642
rect 2732 3056 2786 3642
rect 2786 3056 2788 3642
rect 2888 3056 2890 3642
rect 2890 3056 2944 3642
rect 2944 3056 2946 3642
rect 3046 3056 3048 3642
rect 3048 3056 3102 3642
rect 3102 3056 3104 3642
rect 3204 3056 3206 3642
rect 3206 3056 3260 3642
rect 3260 3056 3262 3642
rect 3340 2372 3540 2572
<< metal3 >>
rect 120 4332 360 4352
rect 120 4132 140 4332
rect 340 4132 360 4332
rect 120 4112 360 4132
rect 178 3382 248 3388
rect 890 3382 950 4352
rect 1750 4346 1930 4352
rect 1750 3958 1756 4346
rect 1924 3958 1930 4346
rect 1750 3952 1930 3958
rect 178 3322 184 3382
rect 242 3322 950 3382
rect 1112 3740 3110 3952
rect 1112 3642 1182 3740
rect 178 3316 248 3322
rect 1112 3056 1118 3642
rect 1176 3056 1182 3642
rect 1112 3050 1182 3056
rect 1270 3642 1340 3648
rect 1270 3056 1276 3642
rect 1334 3056 1340 3642
rect 1270 2958 1340 3056
rect 1428 3642 1498 3740
rect 1428 3056 1434 3642
rect 1492 3056 1498 3642
rect 1428 3050 1498 3056
rect 1586 3642 1656 3648
rect 1586 3056 1592 3642
rect 1650 3056 1656 3642
rect 1586 2958 1656 3056
rect 1744 3642 1814 3740
rect 1744 3056 1750 3642
rect 1808 3056 1814 3642
rect 1744 3050 1814 3056
rect 2092 3642 2162 3740
rect 2092 3056 2098 3642
rect 2156 3056 2162 3642
rect 2092 3050 2162 3056
rect 2250 3642 2320 3648
rect 2250 3056 2256 3642
rect 2314 3056 2320 3642
rect 2250 2958 2320 3056
rect 2408 3642 2478 3740
rect 2408 3056 2414 3642
rect 2472 3056 2478 3642
rect 2408 3050 2478 3056
rect 2566 3642 2636 3648
rect 2566 3056 2572 3642
rect 2630 3056 2636 3642
rect 2566 2958 2636 3056
rect 2724 3642 2794 3740
rect 2724 3056 2730 3642
rect 2788 3056 2794 3642
rect 2724 3050 2794 3056
rect 2882 3642 2952 3648
rect 2882 3056 2888 3642
rect 2946 3056 2952 3642
rect 2882 2958 2952 3056
rect 3040 3642 3110 3740
rect 3040 3056 3046 3642
rect 3104 3056 3110 3642
rect 3040 3050 3110 3056
rect 3198 3642 3268 3648
rect 3198 3056 3204 3642
rect 3262 3056 3268 3642
rect 3198 2958 3268 3056
rect 1270 2752 3268 2958
rect 1750 2746 1930 2752
rect 1750 2358 1756 2746
rect 1924 2358 1930 2746
rect 1750 2352 1930 2358
rect 3320 2572 3560 2592
rect 3320 2372 3340 2572
rect 3540 2372 3560 2572
rect 3320 2352 3560 2372
<< via3 >>
rect 140 4132 340 4332
rect 1756 3958 1924 4346
rect 1756 2358 1924 2746
rect 3340 2372 3540 2572
<< metal4 >>
rect 120 4332 360 4352
rect 120 4132 140 4332
rect 340 4132 360 4332
rect 120 0 360 4132
rect 1750 4346 1930 4352
rect 1750 3958 1756 4346
rect 1924 3958 1930 4346
rect 1750 3952 1930 3958
rect 1750 2746 1930 2752
rect 1750 2358 1756 2746
rect 1924 2358 1930 2746
rect 1750 2352 1930 2358
rect 3320 2572 3560 4352
rect 3320 2372 3340 2572
rect 3540 2372 3560 2572
rect 3320 0 3560 2372
use sky130_fd_pr__nfet_01v8_lvt_F7BGX5  sky130_fd_pr__nfet_01v8_lvt_F7BGX5_0
timestamp 1712309281
transform 1 0 1463 0 1 3350
box -483 -510 483 510
use sky130_fd_pr__nfet_01v8_NRQ53D  sky130_fd_pr__nfet_01v8_NRQ53D_0
timestamp 1712308627
transform 1 0 665 0 1 3732
box -211 -360 211 360
use sky130_fd_pr__nfet_01v8_NRQ53D  sky130_fd_pr__nfet_01v8_NRQ53D_1
timestamp 1712308627
transform 1 0 349 0 1 3732
box -211 -360 211 360
use sky130_fd_pr__pfet_01v8_lvt_3LP7Y6  sky130_fd_pr__pfet_01v8_lvt_3LP7Y6_1
timestamp 1712309281
transform 1 0 2680 0 1 3349
box -720 -519 720 519
use sky130_fd_pr__pfet_01v8_XJBLHL  sky130_fd_pr__pfet_01v8_XJBLHL_0
timestamp 1712317355
transform 1 0 297 0 1 2963
box -263 -369 263 369
use sky130_fd_pr__pfet_01v8_XJBLHL  sky130_fd_pr__pfet_01v8_XJBLHL_1
timestamp 1712317355
transform 1 0 717 0 1 2963
box -263 -369 263 369
<< labels >>
rlabel metal4 120 0 360 4352 1 VGND
port 1 n ground input
rlabel metal4 3320 0 3560 4352 1 VPWR
port 2 n power input
rlabel metal4 1750 3952 1930 4352 1 mod
port 3 n analog bidirectional
rlabel metal4 1750 2352 1930 2752 1 bus
port 4 n analog bidirectional
rlabel metal3 890 4172 950 4352 1 ctrl
port 5 n signal input
<< properties >>
string FIXED_BBOX 0 0 3680 4352
<< end >>
